// initial begin
assign image [0][0]=	0	;
assign image [0][1]=	0	;
assign image [0][2]=	0	;
assign image [0][3]=	0	;
assign image [0][4]=	0	;
assign image [0][5]=	0	;
assign image [0][6]=	0	;
assign image [0][7]=	0	;
assign image [0][8]=	0	;
assign image [0][9]=	0	;
assign image [0][10]=	0	;
assign image [0][11]=	0	;
assign image [0][12]=	0	;
assign image [0][13]=	0	;
assign image [0][14]=	0	;
assign image [0][15]=	0	;
assign image [0][16]=	0	;
assign image [0][17]=	0	;
assign image [0][18]=	0	;
assign image [0][19]=	0	;
assign image [0][20]=	0	;
assign image [0][21]=	0	;
assign image [0][22]=	0	;
assign image [0][23]=	0	;
assign image [0][24]=	0	;
assign image [0][25]=	0	;
assign image [0][26]=	0	;
assign image [0][27]=	0	;
assign image [1][0]=	0	;
assign image [1][1]=	0	;
assign image [1][2]=	0	;
assign image [1][3]=	0	;
assign image [1][4]=	0	;
assign image [1][5]=	0	;
assign image [1][6]=	0	;
assign image [1][7]=	0	;
assign image [1][8]=	0	;
assign image [1][9]=	0	;
assign image [1][10]=	0	;
assign image [1][11]=	0	;
assign image [1][12]=	0	;
assign image [1][13]=	0	;
assign image [1][14]=	0	;
assign image [1][15]=	0	;
assign image [1][16]=	0	;
assign image [1][17]=	0	;
assign image [1][18]=	0	;
assign image [1][19]=	0	;
assign image [1][20]=	0	;
assign image [1][21]=	0	;
assign image [1][22]=	0	;
assign image [1][23]=	0	;
assign image [1][24]=	0	;
assign image [1][25]=	0	;
assign image [1][26]=	0	;
assign image [1][27]=	0	;
assign image [2][0]=	0	;
assign image [2][1]=	0	;
assign image [2][2]=	0	;
assign image [2][3]=	0	;
assign image [2][4]=	0	;
assign image [2][5]=	0	;
assign image [2][6]=	0	;
assign image [2][7]=	0	;
assign image [2][8]=	0	;
assign image [2][9]=	0	;
assign image [2][10]=	0	;
assign image [2][11]=	0	;
assign image [2][12]=	0	;
assign image [2][13]=	0	;
assign image [2][14]=	0	;
assign image [2][15]=	0	;
assign image [2][16]=	0	;
assign image [2][17]=	0	;
assign image [2][18]=	0	;
assign image [2][19]=	0	;
assign image [2][20]=	0	;
assign image [2][21]=	0	;
assign image [2][22]=	0	;
assign image [2][23]=	0	;
assign image [2][24]=	0	;
assign image [2][25]=	0	;
assign image [2][26]=	0	;
assign image [2][27]=	0	;
assign image [3][0]=	0	;
assign image [3][1]=	0	;
assign image [3][2]=	0	;
assign image [3][3]=	0	;
assign image [3][4]=	0	;
assign image [3][5]=	0	;
assign image [3][6]=	0	;
assign image [3][7]=	0	;
assign image [3][8]=	0	;
assign image [3][9]=	0	;
assign image [3][10]=	0	;
assign image [3][11]=	0	;
assign image [3][12]=	0	;
assign image [3][13]=	0	;
assign image [3][14]=	0	;
assign image [3][15]=	0	;
assign image [3][16]=	0	;
assign image [3][17]=	0	;
assign image [3][18]=	0	;
assign image [3][19]=	0	;
assign image [3][20]=	0	;
assign image [3][21]=	0	;
assign image [3][22]=	0	;
assign image [3][23]=	0	;
assign image [3][24]=	0	;
assign image [3][25]=	0	;
assign image [3][26]=	0	;
assign image [3][27]=	0	;
assign image [4][0]=	0	;
assign image [4][1]=	0	;
assign image [4][2]=	0	;
assign image [4][3]=	0	;
assign image [4][4]=	0	;
assign image [4][5]=	0	;
assign image [4][6]=	0	;
assign image [4][7]=	0	;
assign image [4][8]=	0	;
assign image [4][9]=	0	;
assign image [4][10]=	0	;
assign image [4][11]=	0	;
assign image [4][12]=	0	;
assign image [4][13]=	0	;
assign image [4][14]=	0	;
assign image [4][15]=	0	;
assign image [4][16]=	0	;
assign image [4][17]=	0	;
assign image [4][18]=	0	;
assign image [4][19]=	0	;
assign image [4][20]=	0	;
assign image [4][21]=	0	;
assign image [4][22]=	0	;
assign image [4][23]=	0	;
assign image [4][24]=	0	;
assign image [4][25]=	0	;
assign image [4][26]=	0	;
assign image [4][27]=	0	;
assign image [5][0]=	0	;
assign image [5][1]=	0	;
assign image [5][2]=	0	;
assign image [5][3]=	0	;
assign image [5][4]=	0	;
assign image [5][5]=	0	;
assign image [5][6]=	0	;
assign image [5][7]=	0	;
assign image [5][8]=	0	;
assign image [5][9]=	0	;
assign image [5][10]=	0	;
assign image [5][11]=	0	;
assign image [5][12]=	0	;
assign image [5][13]=	0	;
assign image [5][14]=	0	;
assign image [5][15]=	0	;
assign image [5][16]=	0	;
assign image [5][17]=	0	;
assign image [5][18]=	0	;
assign image [5][19]=	0	;
assign image [5][20]=	67	;
assign image [5][21]=	232	;
assign image [5][22]=	39	;
assign image [5][23]=	0	;
assign image [5][24]=	0	;
assign image [5][25]=	0	;
assign image [5][26]=	0	;
assign image [5][27]=	0	;
assign image [6][0]=	0	;
assign image [6][1]=	0	;
assign image [6][2]=	0	;
assign image [6][3]=	0	;
assign image [6][4]=	62	;
assign image [6][5]=	81	;
assign image [6][6]=	0	;
assign image [6][7]=	0	;
assign image [6][8]=	0	;
assign image [6][9]=	0	;
assign image [6][10]=	0	;
assign image [6][11]=	0	;
assign image [6][12]=	0	;
assign image [6][13]=	0	;
assign image [6][14]=	0	;
assign image [6][15]=	0	;
assign image [6][16]=	0	;
assign image [6][17]=	0	;
assign image [6][18]=	0	;
assign image [6][19]=	0	;
assign image [6][20]=	120	;
assign image [6][21]=	180	;
assign image [6][22]=	39	;
assign image [6][23]=	0	;
assign image [6][24]=	0	;
assign image [6][25]=	0	;
assign image [6][26]=	0	;
assign image [6][27]=	0	;
assign image [7][0]=	0	;
assign image [7][1]=	0	;
assign image [7][2]=	0	;
assign image [7][3]=	0	;
assign image [7][4]=	126	;
assign image [7][5]=	163	;
assign image [7][6]=	0	;
assign image [7][7]=	0	;
assign image [7][8]=	0	;
assign image [7][9]=	0	;
assign image [7][10]=	0	;
assign image [7][11]=	0	;
assign image [7][12]=	0	;
assign image [7][13]=	0	;
assign image [7][14]=	0	;
assign image [7][15]=	0	;
assign image [7][16]=	0	;
assign image [7][17]=	0	;
assign image [7][18]=	0	;
assign image [7][19]=	2	;
assign image [7][20]=	153	;
assign image [7][21]=	210	;
assign image [7][22]=	40	;
assign image [7][23]=	0	;
assign image [7][24]=	0	;
assign image [7][25]=	0	;
assign image [7][26]=	0	;
assign image [7][27]=	0	;
assign image [8][0]=	0	;
assign image [8][1]=	0	;
assign image [8][2]=	0	;
assign image [8][3]=	0	;
assign image [8][4]=	220	;
assign image [8][5]=	163	;
assign image [8][6]=	0	;
assign image [8][7]=	0	;
assign image [8][8]=	0	;
assign image [8][9]=	0	;
assign image [8][10]=	0	;
assign image [8][11]=	0	;
assign image [8][12]=	0	;
assign image [8][13]=	0	;
assign image [8][14]=	0	;
assign image [8][15]=	0	;
assign image [8][16]=	0	;
assign image [8][17]=	0	;
assign image [8][18]=	0	;
assign image [8][19]=	27	;
assign image [8][20]=	254	;
assign image [8][21]=	162	;
assign image [8][22]=	0	;
assign image [8][23]=	0	;
assign image [8][24]=	0	;
assign image [8][25]=	0	;
assign image [8][26]=	0	;
assign image [8][27]=	0	;
assign image [9][0]=	0	;
assign image [9][1]=	0	;
assign image [9][2]=	0	;
assign image [9][3]=	0	;
assign image [9][4]=	222	;
assign image [9][5]=	163	;
assign image [9][6]=	0	;
assign image [9][7]=	0	;
assign image [9][8]=	0	;
assign image [9][9]=	0	;
assign image [9][10]=	0	;
assign image [9][11]=	0	;
assign image [9][12]=	0	;
assign image [9][13]=	0	;
assign image [9][14]=	0	;
assign image [9][15]=	0	;
assign image [9][16]=	0	;
assign image [9][17]=	0	;
assign image [9][18]=	0	;
assign image [9][19]=	183	;
assign image [9][20]=	254	;
assign image [9][21]=	125	;
assign image [9][22]=	0	;
assign image [9][23]=	0	;
assign image [9][24]=	0	;
assign image [9][25]=	0	;
assign image [9][26]=	0	;
assign image [9][27]=	0	;
assign image [10][0]=	0	;
assign image [10][1]=	0	;
assign image [10][2]=	0	;
assign image [10][3]=	46	;
assign image [10][4]=	245	;
assign image [10][5]=	163	;
assign image [10][6]=	0	;
assign image [10][7]=	0	;
assign image [10][8]=	0	;
assign image [10][9]=	0	;
assign image [10][10]=	0	;
assign image [10][11]=	0	;
assign image [10][12]=	0	;
assign image [10][13]=	0	;
assign image [10][14]=	0	;
assign image [10][15]=	0	;
assign image [10][16]=	0	;
assign image [10][17]=	0	;
assign image [10][18]=	0	;
assign image [10][19]=	198	;
assign image [10][20]=	254	;
assign image [10][21]=	56	;
assign image [10][22]=	0	;
assign image [10][23]=	0	;
assign image [10][24]=	0	;
assign image [10][25]=	0	;
assign image [10][26]=	0	;
assign image [10][27]=	0	;
assign image [11][0]=	0	;
assign image [11][1]=	0	;
assign image [11][2]=	0	;
assign image [11][3]=	120	;
assign image [11][4]=	254	;
assign image [11][5]=	163	;
assign image [11][6]=	0	;
assign image [11][7]=	0	;
assign image [11][8]=	0	;
assign image [11][9]=	0	;
assign image [11][10]=	0	;
assign image [11][11]=	0	;
assign image [11][12]=	0	;
assign image [11][13]=	0	;
assign image [11][14]=	0	;
assign image [11][15]=	0	;
assign image [11][16]=	0	;
assign image [11][17]=	0	;
assign image [11][18]=	23	;
assign image [11][19]=	231	;
assign image [11][20]=	254	;
assign image [11][21]=	29	;
assign image [11][22]=	0	;
assign image [11][23]=	0	;
assign image [11][24]=	0	;
assign image [11][25]=	0	;
assign image [11][26]=	0	;
assign image [11][27]=	0	;
assign image [12][0]=	0	;
assign image [12][1]=	0	;
assign image [12][2]=	0	;
assign image [12][3]=	159	;
assign image [12][4]=	254	;
assign image [12][5]=	120	;
assign image [12][6]=	0	;
assign image [12][7]=	0	;
assign image [12][8]=	0	;
assign image [12][9]=	0	;
assign image [12][10]=	0	;
assign image [12][11]=	0	;
assign image [12][12]=	0	;
assign image [12][13]=	0	;
assign image [12][14]=	0	;
assign image [12][15]=	0	;
assign image [12][16]=	0	;
assign image [12][17]=	0	;
assign image [12][18]=	163	;
assign image [12][19]=	254	;
assign image [12][20]=	216	;
assign image [12][21]=	16	;
assign image [12][22]=	0	;
assign image [12][23]=	0	;
assign image [12][24]=	0	;
assign image [12][25]=	0	;
assign image [12][26]=	0	;
assign image [12][27]=	0	;
assign image [13][0]=	0	;
assign image [13][1]=	0	;
assign image [13][2]=	0	;
assign image [13][3]=	159	;
assign image [13][4]=	254	;
assign image [13][5]=	67	;
assign image [13][6]=	0	;
assign image [13][7]=	0	;
assign image [13][8]=	0	;
assign image [13][9]=	0	;
assign image [13][10]=	0	;
assign image [13][11]=	0	;
assign image [13][12]=	0	;
assign image [13][13]=	0	;
assign image [13][14]=	0	;
assign image [13][15]=	14	;
assign image [13][16]=	86	;
assign image [13][17]=	178	;
assign image [13][18]=	248	;
assign image [13][19]=	254	;
assign image [13][20]=	91	;
assign image [13][21]=	0	;
assign image [13][22]=	0	;
assign image [13][23]=	0	;
assign image [13][24]=	0	;
assign image [13][25]=	0	;
assign image [13][26]=	0	;
assign image [13][27]=	0	;
assign image [14][0]=	0	;
assign image [14][1]=	0	;
assign image [14][2]=	0	;
assign image [14][3]=	159	;
assign image [14][4]=	254	;
assign image [14][5]=	85	;
assign image [14][6]=	0	;
assign image [14][7]=	0	;
assign image [14][8]=	0	;
assign image [14][9]=	47	;
assign image [14][10]=	49	;
assign image [14][11]=	116	;
assign image [14][12]=	144	;
assign image [14][13]=	150	;
assign image [14][14]=	241	;
assign image [14][15]=	243	;
assign image [14][16]=	234	;
assign image [14][17]=	179	;
assign image [14][18]=	241	;
assign image [14][19]=	252	;
assign image [14][20]=	40	;
assign image [14][21]=	0	;
assign image [14][22]=	0	;
assign image [14][23]=	0	;
assign image [14][24]=	0	;
assign image [14][25]=	0	;
assign image [14][26]=	0	;
assign image [14][27]=	0	;
assign image [15][0]=	0	;
assign image [15][1]=	0	;
assign image [15][2]=	0	;
assign image [15][3]=	150	;
assign image [15][4]=	253	;
assign image [15][5]=	237	;
assign image [15][6]=	207	;
assign image [15][7]=	207	;
assign image [15][8]=	207	;
assign image [15][9]=	253	;
assign image [15][10]=	254	;
assign image [15][11]=	250	;
assign image [15][12]=	240	;
assign image [15][13]=	198	;
assign image [15][14]=	143	;
assign image [15][15]=	91	;
assign image [15][16]=	28	;
assign image [15][17]=	5	;
assign image [15][18]=	233	;
assign image [15][19]=	250	;
assign image [15][20]=	0	;
assign image [15][21]=	0	;
assign image [15][22]=	0	;
assign image [15][23]=	0	;
assign image [15][24]=	0	;
assign image [15][25]=	0	;
assign image [15][26]=	0	;
assign image [15][27]=	0	;
assign image [16][0]=	0	;
assign image [16][1]=	0	;
assign image [16][2]=	0	;
assign image [16][3]=	0	;
assign image [16][4]=	119	;
assign image [16][5]=	177	;
assign image [16][6]=	177	;
assign image [16][7]=	177	;
assign image [16][8]=	177	;
assign image [16][9]=	177	;
assign image [16][10]=	98	;
assign image [16][11]=	56	;
assign image [16][12]=	0	;
assign image [16][13]=	0	;
assign image [16][14]=	0	;
assign image [16][15]=	0	;
assign image [16][16]=	0	;
assign image [16][17]=	102	;
assign image [16][18]=	254	;
assign image [16][19]=	220	;
assign image [16][20]=	0	;
assign image [16][21]=	0	;
assign image [16][22]=	0	;
assign image [16][23]=	0	;
assign image [16][24]=	0	;
assign image [16][25]=	0	;
assign image [16][26]=	0	;
assign image [16][27]=	0	;
assign image [17][0]=	0	;
assign image [17][1]=	0	;
assign image [17][2]=	0	;
assign image [17][3]=	0	;
assign image [17][4]=	0	;
assign image [17][5]=	0	;
assign image [17][6]=	0	;
assign image [17][7]=	0	;
assign image [17][8]=	0	;
assign image [17][9]=	0	;
assign image [17][10]=	0	;
assign image [17][11]=	0	;
assign image [17][12]=	0	;
assign image [17][13]=	0	;
assign image [17][14]=	0	;
assign image [17][15]=	0	;
assign image [17][16]=	0	;
assign image [17][17]=	169	;
assign image [17][18]=	254	;
assign image [17][19]=	137	;
assign image [17][20]=	0	;
assign image [17][21]=	0	;
assign image [17][22]=	0	;
assign image [17][23]=	0	;
assign image [17][24]=	0	;
assign image [17][25]=	0	;
assign image [17][26]=	0	;
assign image [17][27]=	0	;
assign image [18][0]=	0	;
assign image [18][1]=	0	;
assign image [18][2]=	0	;
assign image [18][3]=	0	;
assign image [18][4]=	0	;
assign image [18][5]=	0	;
assign image [18][6]=	0	;
assign image [18][7]=	0	;
assign image [18][8]=	0	;
assign image [18][9]=	0	;
assign image [18][10]=	0	;
assign image [18][11]=	0	;
assign image [18][12]=	0	;
assign image [18][13]=	0	;
assign image [18][14]=	0	;
assign image [18][15]=	0	;
assign image [18][16]=	0	;
assign image [18][17]=	169	;
assign image [18][18]=	254	;
assign image [18][19]=	57	;
assign image [18][20]=	0	;
assign image [18][21]=	0	;
assign image [18][22]=	0	;
assign image [18][23]=	0	;
assign image [18][24]=	0	;
assign image [18][25]=	0	;
assign image [18][26]=	0	;
assign image [18][27]=	0	;
assign image [19][0]=	0	;
assign image [19][1]=	0	;
assign image [19][2]=	0	;
assign image [19][3]=	0	;
assign image [19][4]=	0	;
assign image [19][5]=	0	;
assign image [19][6]=	0	;
assign image [19][7]=	0	;
assign image [19][8]=	0	;
assign image [19][9]=	0	;
assign image [19][10]=	0	;
assign image [19][11]=	0	;
assign image [19][12]=	0	;
assign image [19][13]=	0	;
assign image [19][14]=	0	;
assign image [19][15]=	0	;
assign image [19][16]=	0	;
assign image [19][17]=	169	;
assign image [19][18]=	254	;
assign image [19][19]=	57	;
assign image [19][20]=	0	;
assign image [19][21]=	0	;
assign image [19][22]=	0	;
assign image [19][23]=	0	;
assign image [19][24]=	0	;
assign image [19][25]=	0	;
assign image [19][26]=	0	;
assign image [19][27]=	0	;
assign image [20][0]=	0	;
assign image [20][1]=	0	;
assign image [20][2]=	0	;
assign image [20][3]=	0	;
assign image [20][4]=	0	;
assign image [20][5]=	0	;
assign image [20][6]=	0	;
assign image [20][7]=	0	;
assign image [20][8]=	0	;
assign image [20][9]=	0	;
assign image [20][10]=	0	;
assign image [20][11]=	0	;
assign image [20][12]=	0	;
assign image [20][13]=	0	;
assign image [20][14]=	0	;
assign image [20][15]=	0	;
assign image [20][16]=	0	;
assign image [20][17]=	169	;
assign image [20][18]=	256	;
assign image [20][19]=	94	;
assign image [20][20]=	0	;
assign image [20][21]=	0	;
assign image [20][22]=	0	;
assign image [20][23]=	0	;
assign image [20][24]=	0	;
assign image [20][25]=	0	;
assign image [20][26]=	0	;
assign image [20][27]=	0	;
assign image [21][0]=	0	;
assign image [21][1]=	0	;
assign image [21][2]=	0	;
assign image [21][3]=	0	;
assign image [21][4]=	0	;
assign image [21][5]=	0	;
assign image [21][6]=	0	;
assign image [21][7]=	0	;
assign image [21][8]=	0	;
assign image [21][9]=	0	;
assign image [21][10]=	0	;
assign image [21][11]=	0	;
assign image [21][12]=	0	;
assign image [21][13]=	0	;
assign image [21][14]=	0	;
assign image [21][15]=	0	;
assign image [21][16]=	0	;
assign image [21][17]=	169	;
assign image [21][18]=	254	;
assign image [21][19]=	96	;
assign image [21][20]=	0	;
assign image [21][21]=	0	;
assign image [21][22]=	0	;
assign image [21][23]=	0	;
assign image [21][24]=	0	;
assign image [21][25]=	0	;
assign image [21][26]=	0	;
assign image [21][27]=	0	;
assign image [22][0]=	0	;
assign image [22][1]=	0	;
assign image [22][2]=	0	;
assign image [22][3]=	0	;
assign image [22][4]=	0	;
assign image [22][5]=	0	;
assign image [22][6]=	0	;
assign image [22][7]=	0	;
assign image [22][8]=	0	;
assign image [22][9]=	0	;
assign image [22][10]=	0	;
assign image [22][11]=	0	;
assign image [22][12]=	0	;
assign image [22][13]=	0	;
assign image [22][14]=	0	;
assign image [22][15]=	0	;
assign image [22][16]=	0	;
assign image [22][17]=	169	;
assign image [22][18]=	254	;
assign image [22][19]=	153	;
assign image [22][20]=	0	;
assign image [22][21]=	0	;
assign image [22][22]=	0	;
assign image [22][23]=	0	;
assign image [22][24]=	0	;
assign image [22][25]=	0	;
assign image [22][26]=	0	;
assign image [22][27]=	0	;
assign image [23][0]=	0	;
assign image [23][1]=	0	;
assign image [23][2]=	0	;
assign image [23][3]=	0	;
assign image [23][4]=	0	;
assign image [23][5]=	0	;
assign image [23][6]=	0	;
assign image [23][7]=	0	;
assign image [23][8]=	0	;
assign image [23][9]=	0	;
assign image [23][10]=	0	;
assign image [23][11]=	0	;
assign image [23][12]=	0	;
assign image [23][13]=	0	;
assign image [23][14]=	0	;
assign image [23][15]=	0	;
assign image [23][16]=	0	;
assign image [23][17]=	169	;
assign image [23][18]=	256	;
assign image [23][19]=	153	;
assign image [23][20]=	0	;
assign image [23][21]=	0	;
assign image [23][22]=	0	;
assign image [23][23]=	0	;
assign image [23][24]=	0	;
assign image [23][25]=	0	;
assign image [23][26]=	0	;
assign image [23][27]=	0	;
assign image [24][0]=	0	;
assign image [24][1]=	0	;
assign image [24][2]=	0	;
assign image [24][3]=	0	;
assign image [24][4]=	0	;
assign image [24][5]=	0	;
assign image [24][6]=	0	;
assign image [24][7]=	0	;
assign image [24][8]=	0	;
assign image [24][9]=	0	;
assign image [24][10]=	0	;
assign image [24][11]=	0	;
assign image [24][12]=	0	;
assign image [24][13]=	0	;
assign image [24][14]=	0	;
assign image [24][15]=	0	;
assign image [24][16]=	0	;
assign image [24][17]=	96	;
assign image [24][18]=	254	;
assign image [24][19]=	153	;
assign image [24][20]=	0	;
assign image [24][21]=	0	;
assign image [24][22]=	0	;
assign image [24][23]=	0	;
assign image [24][24]=	0	;
assign image [24][25]=	0	;
assign image [24][26]=	0	;
assign image [24][27]=	0	;
assign image [25][0]=	0	;
assign image [25][1]=	0	;
assign image [25][2]=	0	;
assign image [25][3]=	0	;
assign image [25][4]=	0	;
assign image [25][5]=	0	;
assign image [25][6]=	0	;
assign image [25][7]=	0	;
assign image [25][8]=	0	;
assign image [25][9]=	0	;
assign image [25][10]=	0	;
assign image [25][11]=	0	;
assign image [25][12]=	0	;
assign image [25][13]=	0	;
assign image [25][14]=	0	;
assign image [25][15]=	0	;
assign image [25][16]=	0	;
assign image [25][17]=	0	;
assign image [25][18]=	0	;
assign image [25][19]=	0	;
assign image [25][20]=	0	;
assign image [25][21]=	0	;
assign image [25][22]=	0	;
assign image [25][23]=	0	;
assign image [25][24]=	0	;
assign image [25][25]=	0	;
assign image [25][26]=	0	;
assign image [25][27]=	0	;
assign image [26][0]=	0	;
assign image [26][1]=	0	;
assign image [26][2]=	0	;
assign image [26][3]=	0	;
assign image [26][4]=	0	;
assign image [26][5]=	0	;
assign image [26][6]=	0	;
assign image [26][7]=	0	;
assign image [26][8]=	0	;
assign image [26][9]=	0	;
assign image [26][10]=	0	;
assign image [26][11]=	0	;
assign image [26][12]=	0	;
assign image [26][13]=	0	;
assign image [26][14]=	0	;
assign image [26][15]=	0	;
assign image [26][16]=	0	;
assign image [26][17]=	0	;
assign image [26][18]=	0	;
assign image [26][19]=	0	;
assign image [26][20]=	0	;
assign image [26][21]=	0	;
assign image [26][22]=	0	;
assign image [26][23]=	0	;
assign image [26][24]=	0	;
assign image [26][25]=	0	;
assign image [26][26]=	0	;
assign image [26][27]=	0	;
assign image [27][0]=	0	;
assign image [27][1]=	0	;
assign image [27][2]=	0	;
assign image [27][3]=	0	;
assign image [27][4]=	0	;
assign image [27][5]=	0	;
assign image [27][6]=	0	;
assign image [27][7]=	0	;
assign image [27][8]=	0	;
assign image [27][9]=	0	;
assign image [27][10]=	0	;
assign image [27][11]=	0	;
assign image [27][12]=	0	;
assign image [27][13]=	0	;
assign image [27][14]=	0	;
assign image [27][15]=	0	;
assign image [27][16]=	0	;
assign image [27][17]=	0	;
assign image [27][18]=	0	;
assign image [27][19]=	0	;
assign image [27][20]=	0	;
assign image [27][21]=	0	;
assign image [27][22]=	0	;
assign image [27][23]=	0	;
assign image [27][24]=	0	;
assign image [27][25]=	0	;
assign image [27][26]=	0	;
assign image [27][27]=	0	;


// end