// module kernel_matrix_trained(conv1_kernel,conv2_kernel,conv3_kernel,connect_matrix);
//     parameter bitwidth=32;
//     output reg signed [bitwidth-1:0] conv1_kernel [1:0][4:0][4:0];
// 	output reg signed [bitwidth-1:0] conv2_kernel [1:0][1:0][4:0][4:0];
// 	output reg signed [bitwidth-1:0] conv3_kernel [9:0][1:0][4:0][4:0];
// 	output reg signed [bitwidth-1:0] connect_matrix [9:0][9:0];
//     always@(*) begin
initial begin
conv1_kernel[0][0][0]=	-146	;
conv1_kernel[0][0][1]=	-101	;
conv1_kernel[0][0][2]=	46	;
conv1_kernel[0][0][3]=	-25	;
conv1_kernel[0][0][4]=	53	;
conv1_kernel[0][1][0]=	-180	;
conv1_kernel[0][1][1]=	48	;
conv1_kernel[0][1][2]=	45	;
conv1_kernel[0][1][3]=	47	;
conv1_kernel[0][1][4]=	25	;
conv1_kernel[0][2][0]=	-142	;
conv1_kernel[0][2][1]=	137	;
conv1_kernel[0][2][2]=	76	;
conv1_kernel[0][2][3]=	73	;
conv1_kernel[0][2][4]=	-10	;
conv1_kernel[0][3][0]=	-54	;
conv1_kernel[0][3][1]=	31	;
conv1_kernel[0][3][2]=	63	;
conv1_kernel[0][3][3]=	33	;
conv1_kernel[0][3][4]=	9	;
conv1_kernel[0][4][0]=	-35	;
conv1_kernel[0][4][1]=	68	;
conv1_kernel[0][4][2]=	-13	;
conv1_kernel[0][4][3]=	-28	;
conv1_kernel[0][4][4]=	-71	;
conv1_kernel[1][0][0]=	28	;
conv1_kernel[1][0][1]=	9	;
conv1_kernel[1][0][2]=	14	;
conv1_kernel[1][0][3]=	-24	;
conv1_kernel[1][0][4]=	-32	;
conv1_kernel[1][1][0]=	53	;
conv1_kernel[1][1][1]=	18	;
conv1_kernel[1][1][2]=	-4	;
conv1_kernel[1][1][3]=	1	;
conv1_kernel[1][1][4]=	-8	;
conv1_kernel[1][2][0]=	46	;
conv1_kernel[1][2][1]=	57	;
conv1_kernel[1][2][2]=	4	;
conv1_kernel[1][2][3]=	1	;
conv1_kernel[1][2][4]=	61	;
conv1_kernel[1][3][0]=	-12	;
conv1_kernel[1][3][1]=	84	;
conv1_kernel[1][3][2]=	134	;
conv1_kernel[1][3][3]=	56	;
conv1_kernel[1][3][4]=	13	;
conv1_kernel[1][4][0]=	-1	;
conv1_kernel[1][4][1]=	-11	;
conv1_kernel[1][4][2]=	4	;
conv1_kernel[1][4][3]=	30	;
conv1_kernel[1][4][4]=	31	;
conv2_kernel[0][0][0][0]=	22	;
conv2_kernel[0][0][0][1]=	54	;
conv2_kernel[0][0][0][2]=	69	;
conv2_kernel[0][0][0][3]=	0	;
conv2_kernel[0][0][0][4]=	-6	;
conv2_kernel[0][0][1][0]=	-70	;
conv2_kernel[0][0][1][1]=	50	;
conv2_kernel[0][0][1][2]=	35	;
conv2_kernel[0][0][1][3]=	-23	;
conv2_kernel[0][0][1][4]=	-24	;
conv2_kernel[0][0][2][0]=	16	;
conv2_kernel[0][0][2][1]=	-29	;
conv2_kernel[0][0][2][2]=	-10	;
conv2_kernel[0][0][2][3]=	6	;
conv2_kernel[0][0][2][4]=	45	;
conv2_kernel[0][0][3][0]=	28	;
conv2_kernel[0][0][3][1]=	5	;
conv2_kernel[0][0][3][2]=	-1	;
conv2_kernel[0][0][3][3]=	60	;
conv2_kernel[0][0][3][4]=	22	;
conv2_kernel[0][0][4][0]=	2	;
conv2_kernel[0][0][4][1]=	-60	;
conv2_kernel[0][0][4][2]=	-79	;
conv2_kernel[0][0][4][3]=	-114	;
conv2_kernel[0][0][4][4]=	-17	;
conv2_kernel[0][1][0][0]=	-61	;
conv2_kernel[0][1][0][1]=	-29	;
conv2_kernel[0][1][0][2]=	8	;
conv2_kernel[0][1][0][3]=	32	;
conv2_kernel[0][1][0][4]=	-55	;
conv2_kernel[0][1][1][0]=	-82	;
conv2_kernel[0][1][1][1]=	0	;
conv2_kernel[0][1][1][2]=	6	;
conv2_kernel[0][1][1][3]=	26	;
conv2_kernel[0][1][1][4]=	62	;
conv2_kernel[0][1][2][0]=	63	;
conv2_kernel[0][1][2][1]=	117	;
conv2_kernel[0][1][2][2]=	137	;
conv2_kernel[0][1][2][3]=	158	;
conv2_kernel[0][1][2][4]=	46	;
conv2_kernel[0][1][3][0]=	-36	;
conv2_kernel[0][1][3][1]=	-54	;
conv2_kernel[0][1][3][2]=	-1	;
conv2_kernel[0][1][3][3]=	-60	;
conv2_kernel[0][1][3][4]=	-181	;
conv2_kernel[0][1][4][0]=	-17	;
conv2_kernel[0][1][4][1]=	19	;
conv2_kernel[0][1][4][2]=	-58	;
conv2_kernel[0][1][4][3]=	-90	;
conv2_kernel[0][1][4][4]=	3	;
conv2_kernel[1][0][0][0]=	81	;
conv2_kernel[1][0][0][1]=	56	;
conv2_kernel[1][0][0][2]=	-30	;
conv2_kernel[1][0][0][3]=	-60	;
conv2_kernel[1][0][0][4]=	-24	;
conv2_kernel[1][0][1][0]=	-68	;
conv2_kernel[1][0][1][1]=	-94	;
conv2_kernel[1][0][1][2]=	55	;
conv2_kernel[1][0][1][3]=	-4	;
conv2_kernel[1][0][1][4]=	-58	;
conv2_kernel[1][0][2][0]=	-75	;
conv2_kernel[1][0][2][1]=	-68	;
conv2_kernel[1][0][2][2]=	46	;
conv2_kernel[1][0][2][3]=	49	;
conv2_kernel[1][0][2][4]=	23	;
conv2_kernel[1][0][3][0]=	19	;
conv2_kernel[1][0][3][1]=	-40	;
conv2_kernel[1][0][3][2]=	-123	;
conv2_kernel[1][0][3][3]=	-7	;
conv2_kernel[1][0][3][4]=	8	;
conv2_kernel[1][0][4][0]=	30	;
conv2_kernel[1][0][4][1]=	17	;
conv2_kernel[1][0][4][2]=	12	;
conv2_kernel[1][0][4][3]=	-5	;
conv2_kernel[1][0][4][4]=	7	;
conv2_kernel[1][1][0][0]=	-95	;
conv2_kernel[1][1][0][1]=	-64	;
conv2_kernel[1][1][0][2]=	-83	;
conv2_kernel[1][1][0][3]=	-86	;
conv2_kernel[1][1][0][4]=	-97	;
conv2_kernel[1][1][1][0]=	-23	;
conv2_kernel[1][1][1][1]=	-117	;
conv2_kernel[1][1][1][2]=	21	;
conv2_kernel[1][1][1][3]=	38	;
conv2_kernel[1][1][1][4]=	71	;
conv2_kernel[1][1][2][0]=	248	;
conv2_kernel[1][1][2][1]=	216	;
conv2_kernel[1][1][2][2]=	94	;
conv2_kernel[1][1][2][3]=	10	;
conv2_kernel[1][1][2][4]=	70	;
conv2_kernel[1][1][3][0]=	-99	;
conv2_kernel[1][1][3][1]=	33	;
conv2_kernel[1][1][3][2]=	0	;
conv2_kernel[1][1][3][3]=	29	;
conv2_kernel[1][1][3][4]=	-22	;
conv2_kernel[1][1][4][0]=	-146	;
conv2_kernel[1][1][4][1]=	-26	;
conv2_kernel[1][1][4][2]=	28	;
conv2_kernel[1][1][4][3]=	20	;
conv2_kernel[1][1][4][4]=	-7	;
conv3_kernel[0][0][0][0]=	-131	;
conv3_kernel[0][0][0][1]=	-30	;
conv3_kernel[0][0][0][2]=	38	;
conv3_kernel[0][0][0][3]=	49	;
conv3_kernel[0][0][0][4]=	11	;
conv3_kernel[0][0][1][0]=	-58	;
conv3_kernel[0][0][1][1]=	-6	;
conv3_kernel[0][0][1][2]=	10	;
conv3_kernel[0][0][1][3]=	-13	;
conv3_kernel[0][0][1][4]=	35	;
conv3_kernel[0][0][2][0]=	56	;
conv3_kernel[0][0][2][1]=	35	;
conv3_kernel[0][0][2][2]=	40	;
conv3_kernel[0][0][2][3]=	14	;
conv3_kernel[0][0][2][4]=	2	;
conv3_kernel[0][0][3][0]=	25	;
conv3_kernel[0][0][3][1]=	-9	;
conv3_kernel[0][0][3][2]=	63	;
conv3_kernel[0][0][3][3]=	-45	;
conv3_kernel[0][0][3][4]=	27	;
conv3_kernel[0][0][4][0]=	13	;
conv3_kernel[0][0][4][1]=	-32	;
conv3_kernel[0][0][4][2]=	14	;
conv3_kernel[0][0][4][3]=	4	;
conv3_kernel[0][0][4][4]=	3	;
conv3_kernel[0][1][0][0]=	-38	;
conv3_kernel[0][1][0][1]=	40	;
conv3_kernel[0][1][0][2]=	28	;
conv3_kernel[0][1][0][3]=	-71	;
conv3_kernel[0][1][0][4]=	-35	;
conv3_kernel[0][1][1][0]=	-144	;
conv3_kernel[0][1][1][1]=	12	;
conv3_kernel[0][1][1][2]=	44	;
conv3_kernel[0][1][1][3]=	4	;
conv3_kernel[0][1][1][4]=	-4	;
conv3_kernel[0][1][2][0]=	-96	;
conv3_kernel[0][1][2][1]=	-9	;
conv3_kernel[0][1][2][2]=	55	;
conv3_kernel[0][1][2][3]=	50	;
conv3_kernel[0][1][2][4]=	-94	;
conv3_kernel[0][1][3][0]=	107	;
conv3_kernel[0][1][3][1]=	6	;
conv3_kernel[0][1][3][2]=	-6	;
conv3_kernel[0][1][3][3]=	-33	;
conv3_kernel[0][1][3][4]=	49	;
conv3_kernel[0][1][4][0]=	164	;
conv3_kernel[0][1][4][1]=	-40	;
conv3_kernel[0][1][4][2]=	7	;
conv3_kernel[0][1][4][3]=	26	;
conv3_kernel[0][1][4][4]=	100	;
conv3_kernel[1][0][0][0]=	74	;
conv3_kernel[1][0][0][1]=	38	;
conv3_kernel[1][0][0][2]=	-11	;
conv3_kernel[1][0][0][3]=	-28	;
conv3_kernel[1][0][0][4]=	-165	;
conv3_kernel[1][0][1][0]=	25	;
conv3_kernel[1][0][1][1]=	24	;
conv3_kernel[1][0][1][2]=	-23	;
conv3_kernel[1][0][1][3]=	-8	;
conv3_kernel[1][0][1][4]=	-162	;
conv3_kernel[1][0][2][0]=	-100	;
conv3_kernel[1][0][2][1]=	-22	;
conv3_kernel[1][0][2][2]=	-1	;
conv3_kernel[1][0][2][3]=	5	;
conv3_kernel[1][0][2][4]=	107	;
conv3_kernel[1][0][3][0]=	-50	;
conv3_kernel[1][0][3][1]=	57	;
conv3_kernel[1][0][3][2]=	78	;
conv3_kernel[1][0][3][3]=	-2	;
conv3_kernel[1][0][3][4]=	83	;
conv3_kernel[1][0][4][0]=	78	;
conv3_kernel[1][0][4][1]=	75	;
conv3_kernel[1][0][4][2]=	-16	;
conv3_kernel[1][0][4][3]=	-21	;
conv3_kernel[1][0][4][4]=	-10	;
conv3_kernel[1][1][0][0]=	-52	;
conv3_kernel[1][1][0][1]=	-50	;
conv3_kernel[1][1][0][2]=	-23	;
conv3_kernel[1][1][0][3]=	-13	;
conv3_kernel[1][1][0][4]=	46	;
conv3_kernel[1][1][1][0]=	42	;
conv3_kernel[1][1][1][1]=	-12	;
conv3_kernel[1][1][1][2]=	-40	;
conv3_kernel[1][1][1][3]=	48	;
conv3_kernel[1][1][1][4]=	27	;
conv3_kernel[1][1][2][0]=	50	;
conv3_kernel[1][1][2][1]=	14	;
conv3_kernel[1][1][2][2]=	-29	;
conv3_kernel[1][1][2][3]=	69	;
conv3_kernel[1][1][2][4]=	-33	;
conv3_kernel[1][1][3][0]=	-70	;
conv3_kernel[1][1][3][1]=	52	;
conv3_kernel[1][1][3][2]=	-25	;
conv3_kernel[1][1][3][3]=	-11	;
conv3_kernel[1][1][3][4]=	33	;
conv3_kernel[1][1][4][0]=	-179	;
conv3_kernel[1][1][4][1]=	42	;
conv3_kernel[1][1][4][2]=	28	;
conv3_kernel[1][1][4][3]=	87	;
conv3_kernel[1][1][4][4]=	79	;
conv3_kernel[2][0][0][0]=	60	;
conv3_kernel[2][0][0][1]=	84	;
conv3_kernel[2][0][0][2]=	-32	;
conv3_kernel[2][0][0][3]=	35	;
conv3_kernel[2][0][0][4]=	-74	;
conv3_kernel[2][0][1][0]=	-32	;
conv3_kernel[2][0][1][1]=	28	;
conv3_kernel[2][0][1][2]=	19	;
conv3_kernel[2][0][1][3]=	-6	;
conv3_kernel[2][0][1][4]=	-86	;
conv3_kernel[2][0][2][0]=	15	;
conv3_kernel[2][0][2][1]=	15	;
conv3_kernel[2][0][2][2]=	-22	;
conv3_kernel[2][0][2][3]=	118	;
conv3_kernel[2][0][2][4]=	69	;
conv3_kernel[2][0][3][0]=	18	;
conv3_kernel[2][0][3][1]=	-4	;
conv3_kernel[2][0][3][2]=	4	;
conv3_kernel[2][0][3][3]=	118	;
conv3_kernel[2][0][3][4]=	35	;
conv3_kernel[2][0][4][0]=	-13	;
conv3_kernel[2][0][4][1]=	-43	;
conv3_kernel[2][0][4][2]=	-60	;
conv3_kernel[2][0][4][3]=	-7	;
conv3_kernel[2][0][4][4]=	30	;
conv3_kernel[2][1][0][0]=	-3	;
conv3_kernel[2][1][0][1]=	0	;
conv3_kernel[2][1][0][2]=	16	;
conv3_kernel[2][1][0][3]=	-1	;
conv3_kernel[2][1][0][4]=	30	;
conv3_kernel[2][1][1][0]=	58	;
conv3_kernel[2][1][1][1]=	20	;
conv3_kernel[2][1][1][2]=	22	;
conv3_kernel[2][1][1][3]=	58	;
conv3_kernel[2][1][1][4]=	19	;
conv3_kernel[2][1][2][0]=	-49	;
conv3_kernel[2][1][2][1]=	-12	;
conv3_kernel[2][1][2][2]=	19	;
conv3_kernel[2][1][2][3]=	94	;
conv3_kernel[2][1][2][4]=	-90	;
conv3_kernel[2][1][3][0]=	-14	;
conv3_kernel[2][1][3][1]=	13	;
conv3_kernel[2][1][3][2]=	30	;
conv3_kernel[2][1][3][3]=	-60	;
conv3_kernel[2][1][3][4]=	-69	;
conv3_kernel[2][1][4][0]=	50	;
conv3_kernel[2][1][4][1]=	-32	;
conv3_kernel[2][1][4][2]=	-68	;
conv3_kernel[2][1][4][3]=	-14	;
conv3_kernel[2][1][4][4]=	-2	;
conv3_kernel[3][0][0][0]=	20	;
conv3_kernel[3][0][0][1]=	-32	;
conv3_kernel[3][0][0][2]=	25	;
conv3_kernel[3][0][0][3]=	-27	;
conv3_kernel[3][0][0][4]=	-40	;
conv3_kernel[3][0][1][0]=	43	;
conv3_kernel[3][0][1][1]=	-22	;
conv3_kernel[3][0][1][2]=	-1	;
conv3_kernel[3][0][1][3]=	2	;
conv3_kernel[3][0][1][4]=	69	;
conv3_kernel[3][0][2][0]=	-1	;
conv3_kernel[3][0][2][1]=	-64	;
conv3_kernel[3][0][2][2]=	1	;
conv3_kernel[3][0][2][3]=	51	;
conv3_kernel[3][0][2][4]=	35	;
conv3_kernel[3][0][3][0]=	-39	;
conv3_kernel[3][0][3][1]=	-18	;
conv3_kernel[3][0][3][2]=	33	;
conv3_kernel[3][0][3][3]=	-117	;
conv3_kernel[3][0][3][4]=	-19	;
conv3_kernel[3][0][4][0]=	65	;
conv3_kernel[3][0][4][1]=	39	;
conv3_kernel[3][0][4][2]=	59	;
conv3_kernel[3][0][4][3]=	-13	;
conv3_kernel[3][0][4][4]=	-64	;
conv3_kernel[3][1][0][0]=	33	;
conv3_kernel[3][1][0][1]=	16	;
conv3_kernel[3][1][0][2]=	17	;
conv3_kernel[3][1][0][3]=	-81	;
conv3_kernel[3][1][0][4]=	34	;
conv3_kernel[3][1][1][0]=	-26	;
conv3_kernel[3][1][1][1]=	4	;
conv3_kernel[3][1][1][2]=	31	;
conv3_kernel[3][1][1][3]=	25	;
conv3_kernel[3][1][1][4]=	-13	;
conv3_kernel[3][1][2][0]=	-32	;
conv3_kernel[3][1][2][1]=	0	;
conv3_kernel[3][1][2][2]=	119	;
conv3_kernel[3][1][2][3]=	85	;
conv3_kernel[3][1][2][4]=	58	;
conv3_kernel[3][1][3][0]=	132	;
conv3_kernel[3][1][3][1]=	-16	;
conv3_kernel[3][1][3][2]=	-19	;
conv3_kernel[3][1][3][3]=	38	;
conv3_kernel[3][1][3][4]=	109	;
conv3_kernel[3][1][4][0]=	-242	;
conv3_kernel[3][1][4][1]=	-26	;
conv3_kernel[3][1][4][2]=	23	;
conv3_kernel[3][1][4][3]=	25	;
conv3_kernel[3][1][4][4]=	-23	;
conv3_kernel[4][0][0][0]=	-15	;
conv3_kernel[4][0][0][1]=	64	;
conv3_kernel[4][0][0][2]=	99	;
conv3_kernel[4][0][0][3]=	156	;
conv3_kernel[4][0][0][4]=	99	;
conv3_kernel[4][0][1][0]=	19	;
conv3_kernel[4][0][1][1]=	7	;
conv3_kernel[4][0][1][2]=	11	;
conv3_kernel[4][0][1][3]=	22	;
conv3_kernel[4][0][1][4]=	48	;
conv3_kernel[4][0][2][0]=	-50	;
conv3_kernel[4][0][2][1]=	-15	;
conv3_kernel[4][0][2][2]=	44	;
conv3_kernel[4][0][2][3]=	-71	;
conv3_kernel[4][0][2][4]=	-90	;
conv3_kernel[4][0][3][0]=	-19	;
conv3_kernel[4][0][3][1]=	3	;
conv3_kernel[4][0][3][2]=	73	;
conv3_kernel[4][0][3][3]=	-47	;
conv3_kernel[4][0][3][4]=	-2	;
conv3_kernel[4][0][4][0]=	17	;
conv3_kernel[4][0][4][1]=	-22	;
conv3_kernel[4][0][4][2]=	39	;
conv3_kernel[4][0][4][3]=	11	;
conv3_kernel[4][0][4][4]=	-58	;
conv3_kernel[4][1][0][0]=	43	;
conv3_kernel[4][1][0][1]=	-30	;
conv3_kernel[4][1][0][2]=	-68	;
conv3_kernel[4][1][0][3]=	-150	;
conv3_kernel[4][1][0][4]=	-35	;
conv3_kernel[4][1][1][0]=	-42	;
conv3_kernel[4][1][1][1]=	-27	;
conv3_kernel[4][1][1][2]=	-13	;
conv3_kernel[4][1][1][3]=	28	;
conv3_kernel[4][1][1][4]=	146	;
conv3_kernel[4][1][2][0]=	-74	;
conv3_kernel[4][1][2][1]=	12	;
conv3_kernel[4][1][2][2]=	61	;
conv3_kernel[4][1][2][3]=	100	;
conv3_kernel[4][1][2][4]=	96	;
conv3_kernel[4][1][3][0]=	-7	;
conv3_kernel[4][1][3][1]=	66	;
conv3_kernel[4][1][3][2]=	9	;
conv3_kernel[4][1][3][3]=	35	;
conv3_kernel[4][1][3][4]=	-20	;
conv3_kernel[4][1][4][0]=	-69	;
conv3_kernel[4][1][4][1]=	46	;
conv3_kernel[4][1][4][2]=	25	;
conv3_kernel[4][1][4][3]=	51	;
conv3_kernel[4][1][4][4]=	-5	;
conv3_kernel[5][0][0][0]=	154	;
conv3_kernel[5][0][0][1]=	67	;
conv3_kernel[5][0][0][2]=	46	;
conv3_kernel[5][0][0][3]=	-34	;
conv3_kernel[5][0][0][4]=	-67	;
conv3_kernel[5][0][1][0]=	89	;
conv3_kernel[5][0][1][1]=	23	;
conv3_kernel[5][0][1][2]=	7	;
conv3_kernel[5][0][1][3]=	-7	;
conv3_kernel[5][0][1][4]=	17	;
conv3_kernel[5][0][2][0]=	30	;
conv3_kernel[5][0][2][1]=	-12	;
conv3_kernel[5][0][2][2]=	-18	;
conv3_kernel[5][0][2][3]=	5	;
conv3_kernel[5][0][2][4]=	-45	;
conv3_kernel[5][0][3][0]=	0	;
conv3_kernel[5][0][3][1]=	26	;
conv3_kernel[5][0][3][2]=	-18	;
conv3_kernel[5][0][3][3]=	-6	;
conv3_kernel[5][0][3][4]=	-4	;
conv3_kernel[5][0][4][0]=	6	;
conv3_kernel[5][0][4][1]=	-47	;
conv3_kernel[5][0][4][2]=	-46	;
conv3_kernel[5][0][4][3]=	17	;
conv3_kernel[5][0][4][4]=	-69	;
conv3_kernel[5][1][0][0]=	-88	;
conv3_kernel[5][1][0][1]=	10	;
conv3_kernel[5][1][0][2]=	32	;
conv3_kernel[5][1][0][3]=	-6	;
conv3_kernel[5][1][0][4]=	12	;
conv3_kernel[5][1][1][0]=	-36	;
conv3_kernel[5][1][1][1]=	61	;
conv3_kernel[5][1][1][2]=	23	;
conv3_kernel[5][1][1][3]=	41	;
conv3_kernel[5][1][1][4]=	18	;
conv3_kernel[5][1][2][0]=	121	;
conv3_kernel[5][1][2][1]=	-14	;
conv3_kernel[5][1][2][2]=	3	;
conv3_kernel[5][1][2][3]=	37	;
conv3_kernel[5][1][2][4]=	75	;
conv3_kernel[5][1][3][0]=	193	;
conv3_kernel[5][1][3][1]=	23	;
conv3_kernel[5][1][3][2]=	-26	;
conv3_kernel[5][1][3][3]=	48	;
conv3_kernel[5][1][3][4]=	20	;
conv3_kernel[5][1][4][0]=	168	;
conv3_kernel[5][1][4][1]=	50	;
conv3_kernel[5][1][4][2]=	38	;
conv3_kernel[5][1][4][3]=	4	;
conv3_kernel[5][1][4][4]=	-42	;
conv3_kernel[6][0][0][0]=	-23	;
conv3_kernel[6][0][0][1]=	-93	;
conv3_kernel[6][0][0][2]=	-48	;
conv3_kernel[6][0][0][3]=	11	;
conv3_kernel[6][0][0][4]=	69	;
conv3_kernel[6][0][1][0]=	-31	;
conv3_kernel[6][0][1][1]=	34	;
conv3_kernel[6][0][1][2]=	18	;
conv3_kernel[6][0][1][3]=	18	;
conv3_kernel[6][0][1][4]=	47	;
conv3_kernel[6][0][2][0]=	35	;
conv3_kernel[6][0][2][1]=	-4	;
conv3_kernel[6][0][2][2]=	-27	;
conv3_kernel[6][0][2][3]=	117	;
conv3_kernel[6][0][2][4]=	37	;
conv3_kernel[6][0][3][0]=	-17	;
conv3_kernel[6][0][3][1]=	37	;
conv3_kernel[6][0][3][2]=	-13	;
conv3_kernel[6][0][3][3]=	48	;
conv3_kernel[6][0][3][4]=	75	;
conv3_kernel[6][0][4][0]=	60	;
conv3_kernel[6][0][4][1]=	-23	;
conv3_kernel[6][0][4][2]=	-1	;
conv3_kernel[6][0][4][3]=	18	;
conv3_kernel[6][0][4][4]=	-19	;
conv3_kernel[6][1][0][0]=	87	;
conv3_kernel[6][1][0][1]=	15	;
conv3_kernel[6][1][0][2]=	-62	;
conv3_kernel[6][1][0][3]=	-143	;
conv3_kernel[6][1][0][4]=	-73	;
conv3_kernel[6][1][1][0]=	-41	;
conv3_kernel[6][1][1][1]=	4	;
conv3_kernel[6][1][1][2]=	-13	;
conv3_kernel[6][1][1][3]=	-21	;
conv3_kernel[6][1][1][4]=	-18	;
conv3_kernel[6][1][2][0]=	79	;
conv3_kernel[6][1][2][1]=	27	;
conv3_kernel[6][1][2][2]=	35	;
conv3_kernel[6][1][2][3]=	136	;
conv3_kernel[6][1][2][4]=	20	;
conv3_kernel[6][1][3][0]=	90	;
conv3_kernel[6][1][3][1]=	30	;
conv3_kernel[6][1][3][2]=	19	;
conv3_kernel[6][1][3][3]=	45	;
conv3_kernel[6][1][3][4]=	97	;
conv3_kernel[6][1][4][0]=	-62	;
conv3_kernel[6][1][4][1]=	-31	;
conv3_kernel[6][1][4][2]=	-23	;
conv3_kernel[6][1][4][3]=	-79	;
conv3_kernel[6][1][4][4]=	44	;
conv3_kernel[7][0][0][0]=	-30	;
conv3_kernel[7][0][0][1]=	-1	;
conv3_kernel[7][0][0][2]=	-83	;
conv3_kernel[7][0][0][3]=	-43	;
conv3_kernel[7][0][0][4]=	-8	;
conv3_kernel[7][0][1][0]=	-142	;
conv3_kernel[7][0][1][1]=	9	;
conv3_kernel[7][0][1][2]=	36	;
conv3_kernel[7][0][1][3]=	18	;
conv3_kernel[7][0][1][4]=	8	;
conv3_kernel[7][0][2][0]=	26	;
conv3_kernel[7][0][2][1]=	25	;
conv3_kernel[7][0][2][2]=	17	;
conv3_kernel[7][0][2][3]=	14	;
conv3_kernel[7][0][2][4]=	33	;
conv3_kernel[7][0][3][0]=	49	;
conv3_kernel[7][0][3][1]=	6	;
conv3_kernel[7][0][3][2]=	-4	;
conv3_kernel[7][0][3][3]=	-46	;
conv3_kernel[7][0][3][4]=	-125	;
conv3_kernel[7][0][4][0]=	-5	;
conv3_kernel[7][0][4][1]=	5	;
conv3_kernel[7][0][4][2]=	-29	;
conv3_kernel[7][0][4][3]=	13	;
conv3_kernel[7][0][4][4]=	67	;
conv3_kernel[7][1][0][0]=	19	;
conv3_kernel[7][1][0][1]=	81	;
conv3_kernel[7][1][0][2]=	10	;
conv3_kernel[7][1][0][3]=	3	;
conv3_kernel[7][1][0][4]=	70	;
conv3_kernel[7][1][1][0]=	78	;
conv3_kernel[7][1][1][1]=	10	;
conv3_kernel[7][1][1][2]=	17	;
conv3_kernel[7][1][1][3]=	18	;
conv3_kernel[7][1][1][4]=	29	;
conv3_kernel[7][1][2][0]=	-75	;
conv3_kernel[7][1][2][1]=	-54	;
conv3_kernel[7][1][2][2]=	68	;
conv3_kernel[7][1][2][3]=	111	;
conv3_kernel[7][1][2][4]=	-13	;
conv3_kernel[7][1][3][0]=	-46	;
conv3_kernel[7][1][3][1]=	48	;
conv3_kernel[7][1][3][2]=	71	;
conv3_kernel[7][1][3][3]=	43	;
conv3_kernel[7][1][3][4]=	-85	;
conv3_kernel[7][1][4][0]=	73	;
conv3_kernel[7][1][4][1]=	40	;
conv3_kernel[7][1][4][2]=	54	;
conv3_kernel[7][1][4][3]=	-20	;
conv3_kernel[7][1][4][4]=	-139	;
conv3_kernel[8][0][0][0]=	-153	;
conv3_kernel[8][0][0][1]=	-59	;
conv3_kernel[8][0][0][2]=	30	;
conv3_kernel[8][0][0][3]=	-7	;
conv3_kernel[8][0][0][4]=	44	;
conv3_kernel[8][0][1][0]=	-232	;
conv3_kernel[8][0][1][1]=	5	;
conv3_kernel[8][0][1][2]=	4	;
conv3_kernel[8][0][1][3]=	10	;
conv3_kernel[8][0][1][4]=	-16	;
conv3_kernel[8][0][2][0]=	45	;
conv3_kernel[8][0][2][1]=	-36	;
conv3_kernel[8][0][2][2]=	32	;
conv3_kernel[8][0][2][3]=	26	;
conv3_kernel[8][0][2][4]=	81	;
conv3_kernel[8][0][3][0]=	-5	;
conv3_kernel[8][0][3][1]=	-6	;
conv3_kernel[8][0][3][2]=	19	;
conv3_kernel[8][0][3][3]=	-31	;
conv3_kernel[8][0][3][4]=	-6	;
conv3_kernel[8][0][4][0]=	35	;
conv3_kernel[8][0][4][1]=	14	;
conv3_kernel[8][0][4][2]=	-4	;
conv3_kernel[8][0][4][3]=	16	;
conv3_kernel[8][0][4][4]=	-10	;
conv3_kernel[8][1][0][0]=	115	;
conv3_kernel[8][1][0][1]=	81	;
conv3_kernel[8][1][0][2]=	6	;
conv3_kernel[8][1][0][3]=	-13	;
conv3_kernel[8][1][0][4]=	61	;
conv3_kernel[8][1][1][0]=	51	;
conv3_kernel[8][1][1][1]=	13	;
conv3_kernel[8][1][1][2]=	20	;
conv3_kernel[8][1][1][3]=	54	;
conv3_kernel[8][1][1][4]=	63	;
conv3_kernel[8][1][2][0]=	12	;
conv3_kernel[8][1][2][1]=	-66	;
conv3_kernel[8][1][2][2]=	-80	;
conv3_kernel[8][1][2][3]=	-31	;
conv3_kernel[8][1][2][4]=	-64	;
conv3_kernel[8][1][3][0]=	-35	;
conv3_kernel[8][1][3][1]=	-28	;
conv3_kernel[8][1][3][2]=	-32	;
conv3_kernel[8][1][3][3]=	-1	;
conv3_kernel[8][1][3][4]=	-54	;
conv3_kernel[8][1][4][0]=	-152	;
conv3_kernel[8][1][4][1]=	19	;
conv3_kernel[8][1][4][2]=	18	;
conv3_kernel[8][1][4][3]=	21	;
conv3_kernel[8][1][4][4]=	-120	;
conv3_kernel[9][0][0][0]=	85	;
conv3_kernel[9][0][0][1]=	-56	;
conv3_kernel[9][0][0][2]=	-57	;
conv3_kernel[9][0][0][3]=	-99	;
conv3_kernel[9][0][0][4]=	-47	;
conv3_kernel[9][0][1][0]=	81	;
conv3_kernel[9][0][1][1]=	-35	;
conv3_kernel[9][0][1][2]=	34	;
conv3_kernel[9][0][1][3]=	36	;
conv3_kernel[9][0][1][4]=	17	;
conv3_kernel[9][0][2][0]=	-6	;
conv3_kernel[9][0][2][1]=	-28	;
conv3_kernel[9][0][2][2]=	140	;
conv3_kernel[9][0][2][3]=	82	;
conv3_kernel[9][0][2][4]=	1	;
conv3_kernel[9][0][3][0]=	-37	;
conv3_kernel[9][0][3][1]=	-31	;
conv3_kernel[9][0][3][2]=	84	;
conv3_kernel[9][0][3][3]=	-60	;
conv3_kernel[9][0][3][4]=	2	;
conv3_kernel[9][0][4][0]=	7	;
conv3_kernel[9][0][4][1]=	-76	;
conv3_kernel[9][0][4][2]=	87	;
conv3_kernel[9][0][4][3]=	48	;
conv3_kernel[9][0][4][4]=	-45	;
conv3_kernel[9][1][0][0]=	-15	;
conv3_kernel[9][1][0][1]=	26	;
conv3_kernel[9][1][0][2]=	89	;
conv3_kernel[9][1][0][3]=	-73	;
conv3_kernel[9][1][0][4]=	-17	;
conv3_kernel[9][1][1][0]=	-9	;
conv3_kernel[9][1][1][1]=	-25	;
conv3_kernel[9][1][1][2]=	23	;
conv3_kernel[9][1][1][3]=	-51	;
conv3_kernel[9][1][1][4]=	-69	;
conv3_kernel[9][1][2][0]=	-5	;
conv3_kernel[9][1][2][1]=	-24	;
conv3_kernel[9][1][2][2]=	57	;
conv3_kernel[9][1][2][3]=	-7	;
conv3_kernel[9][1][2][4]=	-2	;
conv3_kernel[9][1][3][0]=	34	;
conv3_kernel[9][1][3][1]=	13	;
conv3_kernel[9][1][3][2]=	9	;
conv3_kernel[9][1][3][3]=	8	;
conv3_kernel[9][1][3][4]=	6	;
conv3_kernel[9][1][4][0]=	29	;
conv3_kernel[9][1][4][1]=	53	;
conv3_kernel[9][1][4][2]=	2	;
conv3_kernel[9][1][4][3]=	-7	;
conv3_kernel[9][1][4][4]=	-26	;
connect_matrix [0][0]=	-87	;
connect_matrix [0][1]=	98	;
connect_matrix [0][2]=	-13	;
connect_matrix [0][3]=	-78	;
connect_matrix [0][4]=	13	;
connect_matrix [0][5]=	-15	;
connect_matrix [0][6]=	-5	;
connect_matrix [0][7]=	-4	;
connect_matrix [0][8]=	51	;
connect_matrix [0][9]=	-48	;
connect_matrix [1][0]=	107	;
connect_matrix [1][1]=	-35	;
connect_matrix [1][2]=	-101	;
connect_matrix [1][3]=	-78	;
connect_matrix [1][4]=	0	;
connect_matrix [1][5]=	38	;
connect_matrix [1][6]=	40	;
connect_matrix [1][7]=	-188	;
connect_matrix [1][8]=	99	;
connect_matrix [1][9]=	147	;
connect_matrix [2][0]=	41	;
connect_matrix [2][1]=	85	;
connect_matrix [2][2]=	-4	;
connect_matrix [2][3]=	37	;
connect_matrix [2][4]=	-91	;
connect_matrix [2][5]=	49	;
connect_matrix [2][6]=	11	;
connect_matrix [2][7]=	-44	;
connect_matrix [2][8]=	-113	;
connect_matrix [2][9]=	-5	;
connect_matrix [3][0]=	-27	;
connect_matrix [3][1]=	-3	;
connect_matrix [3][2]=	-65	;
connect_matrix [3][3]=	-1	;
connect_matrix [3][4]=	-17	;
connect_matrix [3][5]=	95	;
connect_matrix [3][6]=	-26	;
connect_matrix [3][7]=	44	;
connect_matrix [3][8]=	-91	;
connect_matrix [3][9]=	45	;
connect_matrix [4][0]=	0	;
connect_matrix [4][1]=	-37	;
connect_matrix [4][2]=	-11	;
connect_matrix [4][3]=	-33	;
connect_matrix [4][4]=	-67	;
connect_matrix [4][5]=	-93	;
connect_matrix [4][6]=	128	;
connect_matrix [4][7]=	56	;
connect_matrix [4][8]=	-39	;
connect_matrix [4][9]=	46	;
connect_matrix [5][0]=	36	;
connect_matrix [5][1]=	-64	;
connect_matrix [5][2]=	-68	;
connect_matrix [5][3]=	-25	;
connect_matrix [5][4]=	85	;
connect_matrix [5][5]=	49	;
connect_matrix [5][6]=	-15	;
connect_matrix [5][7]=	40	;
connect_matrix [5][8]=	-13	;
connect_matrix [5][9]=	-75	;
connect_matrix [6][0]=	-105	;
connect_matrix [6][1]=	52	;
connect_matrix [6][2]=	41	;
connect_matrix [6][3]=	19	;
connect_matrix [6][4]=	123	;
connect_matrix [6][5]=	-182	;
connect_matrix [6][6]=	26	;
connect_matrix [6][7]=	-27	;
connect_matrix [6][8]=	-29	;
connect_matrix [6][9]=	-31	;
connect_matrix [7][0]=	-63	;
connect_matrix [7][1]=	-87	;
connect_matrix [7][2]=	108	;
connect_matrix [7][3]=	39	;
connect_matrix [7][4]=	-10	;
connect_matrix [7][5]=	56	;
connect_matrix [7][6]=	-1	;
connect_matrix [7][7]=	-78	;
connect_matrix [7][8]=	55	;
connect_matrix [7][9]=	33	;
connect_matrix [8][0]=	14	;
connect_matrix [8][1]=	-4	;
connect_matrix [8][2]=	5	;
connect_matrix [8][3]=	115	;
connect_matrix [8][4]=	-27	;
connect_matrix [8][5]=	-19	;
connect_matrix [8][6]=	-57	;
connect_matrix [8][7]=	23	;
connect_matrix [8][8]=	22	;
connect_matrix [8][9]=	-18	;
connect_matrix [9][0]=	54	;
connect_matrix [9][1]=	-14	;
connect_matrix [9][2]=	75	;
connect_matrix [9][3]=	-40	;
connect_matrix [9][4]=	-23	;
connect_matrix [9][5]=	-47	;
connect_matrix [9][6]=	-71	;
connect_matrix [9][7]=	85	;
connect_matrix [9][8]=	-63	;
connect_matrix [9][9]=	34	;




end
//     end
// endmodule