// module kernel_matrix_trained(conv1_kernel,conv2_kernel,conv3_kernel,connect_matrix);
//     parameter bitwidth=32;
//     output reg signed [bitwidth-1:0] conv1_kernel [1:0][4:0][4:0];
// 	output reg signed [bitwidth-1:0] conv2_kernel [1:0][1:0][4:0][4:0];
// 	output reg signed [bitwidth-1:0] conv3_kernel [9:0][1:0][4:0][4:0];
// 	output reg signed [bitwidth-1:0] connect_matrix [9:0][9:0];
//     always@(*) begin
// initial begin
assign conv1_kernel[0][0][0]=	-73	;
assign conv1_kernel[0][0][1]=	-51	;
assign conv1_kernel[0][0][2]=	23	;
assign conv1_kernel[0][0][3]=	-12	;
assign conv1_kernel[0][0][4]=	27	;
assign conv1_kernel[0][1][0]=	-90	;
assign conv1_kernel[0][1][1]=	24	;
assign conv1_kernel[0][1][2]=	23	;
assign conv1_kernel[0][1][3]=	23	;
assign conv1_kernel[0][1][4]=	13	;
assign conv1_kernel[0][2][0]=	-71	;
assign conv1_kernel[0][2][1]=	69	;
assign conv1_kernel[0][2][2]=	38	;
assign conv1_kernel[0][2][3]=	37	;
assign conv1_kernel[0][2][4]=	-5	;
assign conv1_kernel[0][3][0]=	-27	;
assign conv1_kernel[0][3][1]=	15	;
assign conv1_kernel[0][3][2]=	32	;
assign conv1_kernel[0][3][3]=	17	;
assign conv1_kernel[0][3][4]=	4	;
assign conv1_kernel[0][4][0]=	-18	;
assign conv1_kernel[0][4][1]=	34	;
assign conv1_kernel[0][4][2]=	-6	;
assign conv1_kernel[0][4][3]=	-14	;
assign conv1_kernel[0][4][4]=	-35	;
assign conv1_kernel[1][0][0]=	14	;
assign conv1_kernel[1][0][1]=	4	;
assign conv1_kernel[1][0][2]=	7	;
assign conv1_kernel[1][0][3]=	-12	;
assign conv1_kernel[1][0][4]=	-16	;
assign conv1_kernel[1][1][0]=	26	;
assign conv1_kernel[1][1][1]=	9	;
assign conv1_kernel[1][1][2]=	-2	;
assign conv1_kernel[1][1][3]=	1	;
assign conv1_kernel[1][1][4]=	-4	;
assign conv1_kernel[1][2][0]=	23	;
assign conv1_kernel[1][2][1]=	28	;
assign conv1_kernel[1][2][2]=	2	;
assign conv1_kernel[1][2][3]=	0	;
assign conv1_kernel[1][2][4]=	30	;
assign conv1_kernel[1][3][0]=	-6	;
assign conv1_kernel[1][3][1]=	42	;
assign conv1_kernel[1][3][2]=	67	;
assign conv1_kernel[1][3][3]=	28	;
assign conv1_kernel[1][3][4]=	6	;
assign conv1_kernel[1][4][0]=	0	;
assign conv1_kernel[1][4][1]=	-6	;
assign conv1_kernel[1][4][2]=	2	;
assign conv1_kernel[1][4][3]=	15	;
assign conv1_kernel[1][4][4]=	15	;
assign conv2_kernel[0][0][0][0]=	11	;
assign conv2_kernel[0][0][0][1]=	27	;
assign conv2_kernel[0][0][0][2]=	34	;
assign conv2_kernel[0][0][0][3]=	0	;
assign conv2_kernel[0][0][0][4]=	-3	;
assign conv2_kernel[0][0][1][0]=	-35	;
assign conv2_kernel[0][0][1][1]=	25	;
assign conv2_kernel[0][0][1][2]=	18	;
assign conv2_kernel[0][0][1][3]=	-11	;
assign conv2_kernel[0][0][1][4]=	-12	;
assign conv2_kernel[0][0][2][0]=	8	;
assign conv2_kernel[0][0][2][1]=	-14	;
assign conv2_kernel[0][0][2][2]=	-5	;
assign conv2_kernel[0][0][2][3]=	3	;
assign conv2_kernel[0][0][2][4]=	22	;
assign conv2_kernel[0][0][3][0]=	14	;
assign conv2_kernel[0][0][3][1]=	2	;
assign conv2_kernel[0][0][3][2]=	-1	;
assign conv2_kernel[0][0][3][3]=	30	;
assign conv2_kernel[0][0][3][4]=	11	;
assign conv2_kernel[0][0][4][0]=	1	;
assign conv2_kernel[0][0][4][1]=	-30	;
assign conv2_kernel[0][0][4][2]=	-39	;
assign conv2_kernel[0][0][4][3]=	-57	;
assign conv2_kernel[0][0][4][4]=	-8	;
assign conv2_kernel[0][1][0][0]=	-30	;
assign conv2_kernel[0][1][0][1]=	-14	;
assign conv2_kernel[0][1][0][2]=	4	;
assign conv2_kernel[0][1][0][3]=	16	;
assign conv2_kernel[0][1][0][4]=	-27	;
assign conv2_kernel[0][1][1][0]=	-41	;
assign conv2_kernel[0][1][1][1]=	0	;
assign conv2_kernel[0][1][1][2]=	3	;
assign conv2_kernel[0][1][1][3]=	13	;
assign conv2_kernel[0][1][1][4]=	31	;
assign conv2_kernel[0][1][2][0]=	32	;
assign conv2_kernel[0][1][2][1]=	58	;
assign conv2_kernel[0][1][2][2]=	69	;
assign conv2_kernel[0][1][2][3]=	79	;
assign conv2_kernel[0][1][2][4]=	23	;
assign conv2_kernel[0][1][3][0]=	-18	;
assign conv2_kernel[0][1][3][1]=	-27	;
assign conv2_kernel[0][1][3][2]=	-1	;
assign conv2_kernel[0][1][3][3]=	-30	;
assign conv2_kernel[0][1][3][4]=	-91	;
assign conv2_kernel[0][1][4][0]=	-9	;
assign conv2_kernel[0][1][4][1]=	10	;
assign conv2_kernel[0][1][4][2]=	-29	;
assign conv2_kernel[0][1][4][3]=	-45	;
assign conv2_kernel[0][1][4][4]=	1	;
assign conv2_kernel[1][0][0][0]=	41	;
assign conv2_kernel[1][0][0][1]=	28	;
assign conv2_kernel[1][0][0][2]=	-15	;
assign conv2_kernel[1][0][0][3]=	-30	;
assign conv2_kernel[1][0][0][4]=	-12	;
assign conv2_kernel[1][0][1][0]=	-34	;
assign conv2_kernel[1][0][1][1]=	-47	;
assign conv2_kernel[1][0][1][2]=	28	;
assign conv2_kernel[1][0][1][3]=	-2	;
assign conv2_kernel[1][0][1][4]=	-29	;
assign conv2_kernel[1][0][2][0]=	-37	;
assign conv2_kernel[1][0][2][1]=	-34	;
assign conv2_kernel[1][0][2][2]=	23	;
assign conv2_kernel[1][0][2][3]=	24	;
assign conv2_kernel[1][0][2][4]=	12	;
assign conv2_kernel[1][0][3][0]=	10	;
assign conv2_kernel[1][0][3][1]=	-20	;
assign conv2_kernel[1][0][3][2]=	-62	;
assign conv2_kernel[1][0][3][3]=	-3	;
assign conv2_kernel[1][0][3][4]=	4	;
assign conv2_kernel[1][0][4][0]=	15	;
assign conv2_kernel[1][0][4][1]=	8	;
assign conv2_kernel[1][0][4][2]=	6	;
assign conv2_kernel[1][0][4][3]=	-3	;
assign conv2_kernel[1][0][4][4]=	4	;
assign conv2_kernel[1][1][0][0]=	-48	;
assign conv2_kernel[1][1][0][1]=	-32	;
assign conv2_kernel[1][1][0][2]=	-41	;
assign conv2_kernel[1][1][0][3]=	-43	;
assign conv2_kernel[1][1][0][4]=	-48	;
assign conv2_kernel[1][1][1][0]=	-12	;
assign conv2_kernel[1][1][1][1]=	-59	;
assign conv2_kernel[1][1][1][2]=	10	;
assign conv2_kernel[1][1][1][3]=	19	;
assign conv2_kernel[1][1][1][4]=	36	;
assign conv2_kernel[1][1][2][0]=	124	;
assign conv2_kernel[1][1][2][1]=	108	;
assign conv2_kernel[1][1][2][2]=	47	;
assign conv2_kernel[1][1][2][3]=	5	;
assign conv2_kernel[1][1][2][4]=	35	;
assign conv2_kernel[1][1][3][0]=	-50	;
assign conv2_kernel[1][1][3][1]=	16	;
assign conv2_kernel[1][1][3][2]=	0	;
assign conv2_kernel[1][1][3][3]=	15	;
assign conv2_kernel[1][1][3][4]=	-11	;
assign conv2_kernel[1][1][4][0]=	-73	;
assign conv2_kernel[1][1][4][1]=	-13	;
assign conv2_kernel[1][1][4][2]=	14	;
assign conv2_kernel[1][1][4][3]=	10	;
assign conv2_kernel[1][1][4][4]=	-3	;
assign conv3_kernel[0][0][0][0]=	-65	;
assign conv3_kernel[0][0][0][1]=	-15	;
assign conv3_kernel[0][0][0][2]=	19	;
assign conv3_kernel[0][0][0][3]=	24	;
assign conv3_kernel[0][0][0][4]=	5	;
assign conv3_kernel[0][0][1][0]=	-29	;
assign conv3_kernel[0][0][1][1]=	-3	;
assign conv3_kernel[0][0][1][2]=	5	;
assign conv3_kernel[0][0][1][3]=	-7	;
assign conv3_kernel[0][0][1][4]=	17	;
assign conv3_kernel[0][0][2][0]=	28	;
assign conv3_kernel[0][0][2][1]=	17	;
assign conv3_kernel[0][0][2][2]=	20	;
assign conv3_kernel[0][0][2][3]=	7	;
assign conv3_kernel[0][0][2][4]=	1	;
assign conv3_kernel[0][0][3][0]=	12	;
assign conv3_kernel[0][0][3][1]=	-5	;
assign conv3_kernel[0][0][3][2]=	32	;
assign conv3_kernel[0][0][3][3]=	-23	;
assign conv3_kernel[0][0][3][4]=	13	;
assign conv3_kernel[0][0][4][0]=	6	;
assign conv3_kernel[0][0][4][1]=	-16	;
assign conv3_kernel[0][0][4][2]=	7	;
assign conv3_kernel[0][0][4][3]=	2	;
assign conv3_kernel[0][0][4][4]=	1	;
assign conv3_kernel[0][1][0][0]=	-19	;
assign conv3_kernel[0][1][0][1]=	20	;
assign conv3_kernel[0][1][0][2]=	14	;
assign conv3_kernel[0][1][0][3]=	-36	;
assign conv3_kernel[0][1][0][4]=	-17	;
assign conv3_kernel[0][1][1][0]=	-72	;
assign conv3_kernel[0][1][1][1]=	6	;
assign conv3_kernel[0][1][1][2]=	22	;
assign conv3_kernel[0][1][1][3]=	2	;
assign conv3_kernel[0][1][1][4]=	-2	;
assign conv3_kernel[0][1][2][0]=	-48	;
assign conv3_kernel[0][1][2][1]=	-4	;
assign conv3_kernel[0][1][2][2]=	27	;
assign conv3_kernel[0][1][2][3]=	25	;
assign conv3_kernel[0][1][2][4]=	-47	;
assign conv3_kernel[0][1][3][0]=	53	;
assign conv3_kernel[0][1][3][1]=	3	;
assign conv3_kernel[0][1][3][2]=	-3	;
assign conv3_kernel[0][1][3][3]=	-17	;
assign conv3_kernel[0][1][3][4]=	25	;
assign conv3_kernel[0][1][4][0]=	82	;
assign conv3_kernel[0][1][4][1]=	-20	;
assign conv3_kernel[0][1][4][2]=	4	;
assign conv3_kernel[0][1][4][3]=	13	;
assign conv3_kernel[0][1][4][4]=	50	;
assign conv3_kernel[1][0][0][0]=	37	;
assign conv3_kernel[1][0][0][1]=	19	;
assign conv3_kernel[1][0][0][2]=	-5	;
assign conv3_kernel[1][0][0][3]=	-14	;
assign conv3_kernel[1][0][0][4]=	-83	;
assign conv3_kernel[1][0][1][0]=	12	;
assign conv3_kernel[1][0][1][1]=	12	;
assign conv3_kernel[1][0][1][2]=	-12	;
assign conv3_kernel[1][0][1][3]=	-4	;
assign conv3_kernel[1][0][1][4]=	-81	;
assign conv3_kernel[1][0][2][0]=	-50	;
assign conv3_kernel[1][0][2][1]=	-11	;
assign conv3_kernel[1][0][2][2]=	-1	;
assign conv3_kernel[1][0][2][3]=	2	;
assign conv3_kernel[1][0][2][4]=	54	;
assign conv3_kernel[1][0][3][0]=	-25	;
assign conv3_kernel[1][0][3][1]=	28	;
assign conv3_kernel[1][0][3][2]=	39	;
assign conv3_kernel[1][0][3][3]=	-1	;
assign conv3_kernel[1][0][3][4]=	41	;
assign conv3_kernel[1][0][4][0]=	39	;
assign conv3_kernel[1][0][4][1]=	37	;
assign conv3_kernel[1][0][4][2]=	-8	;
assign conv3_kernel[1][0][4][3]=	-11	;
assign conv3_kernel[1][0][4][4]=	-5	;
assign conv3_kernel[1][1][0][0]=	-26	;
assign conv3_kernel[1][1][0][1]=	-25	;
assign conv3_kernel[1][1][0][2]=	-12	;
assign conv3_kernel[1][1][0][3]=	-7	;
assign conv3_kernel[1][1][0][4]=	23	;
assign conv3_kernel[1][1][1][0]=	21	;
assign conv3_kernel[1][1][1][1]=	-6	;
assign conv3_kernel[1][1][1][2]=	-20	;
assign conv3_kernel[1][1][1][3]=	24	;
assign conv3_kernel[1][1][1][4]=	13	;
assign conv3_kernel[1][1][2][0]=	25	;
assign conv3_kernel[1][1][2][1]=	7	;
assign conv3_kernel[1][1][2][2]=	-14	;
assign conv3_kernel[1][1][2][3]=	34	;
assign conv3_kernel[1][1][2][4]=	-16	;
assign conv3_kernel[1][1][3][0]=	-35	;
assign conv3_kernel[1][1][3][1]=	26	;
assign conv3_kernel[1][1][3][2]=	-12	;
assign conv3_kernel[1][1][3][3]=	-6	;
assign conv3_kernel[1][1][3][4]=	16	;
assign conv3_kernel[1][1][4][0]=	-90	;
assign conv3_kernel[1][1][4][1]=	21	;
assign conv3_kernel[1][1][4][2]=	14	;
assign conv3_kernel[1][1][4][3]=	43	;
assign conv3_kernel[1][1][4][4]=	39	;
assign conv3_kernel[2][0][0][0]=	30	;
assign conv3_kernel[2][0][0][1]=	42	;
assign conv3_kernel[2][0][0][2]=	-16	;
assign conv3_kernel[2][0][0][3]=	18	;
assign conv3_kernel[2][0][0][4]=	-37	;
assign conv3_kernel[2][0][1][0]=	-16	;
assign conv3_kernel[2][0][1][1]=	14	;
assign conv3_kernel[2][0][1][2]=	10	;
assign conv3_kernel[2][0][1][3]=	-3	;
assign conv3_kernel[2][0][1][4]=	-43	;
assign conv3_kernel[2][0][2][0]=	7	;
assign conv3_kernel[2][0][2][1]=	7	;
assign conv3_kernel[2][0][2][2]=	-11	;
assign conv3_kernel[2][0][2][3]=	59	;
assign conv3_kernel[2][0][2][4]=	35	;
assign conv3_kernel[2][0][3][0]=	9	;
assign conv3_kernel[2][0][3][1]=	-2	;
assign conv3_kernel[2][0][3][2]=	2	;
assign conv3_kernel[2][0][3][3]=	59	;
assign conv3_kernel[2][0][3][4]=	17	;
assign conv3_kernel[2][0][4][0]=	-6	;
assign conv3_kernel[2][0][4][1]=	-22	;
assign conv3_kernel[2][0][4][2]=	-30	;
assign conv3_kernel[2][0][4][3]=	-4	;
assign conv3_kernel[2][0][4][4]=	15	;
assign conv3_kernel[2][1][0][0]=	-2	;
assign conv3_kernel[2][1][0][1]=	0	;
assign conv3_kernel[2][1][0][2]=	8	;
assign conv3_kernel[2][1][0][3]=	0	;
assign conv3_kernel[2][1][0][4]=	15	;
assign conv3_kernel[2][1][1][0]=	29	;
assign conv3_kernel[2][1][1][1]=	10	;
assign conv3_kernel[2][1][1][2]=	11	;
assign conv3_kernel[2][1][1][3]=	29	;
assign conv3_kernel[2][1][1][4]=	10	;
assign conv3_kernel[2][1][2][0]=	-24	;
assign conv3_kernel[2][1][2][1]=	-6	;
assign conv3_kernel[2][1][2][2]=	9	;
assign conv3_kernel[2][1][2][3]=	47	;
assign conv3_kernel[2][1][2][4]=	-45	;
assign conv3_kernel[2][1][3][0]=	-7	;
assign conv3_kernel[2][1][3][1]=	7	;
assign conv3_kernel[2][1][3][2]=	15	;
assign conv3_kernel[2][1][3][3]=	-30	;
assign conv3_kernel[2][1][3][4]=	-35	;
assign conv3_kernel[2][1][4][0]=	25	;
assign conv3_kernel[2][1][4][1]=	-16	;
assign conv3_kernel[2][1][4][2]=	-34	;
assign conv3_kernel[2][1][4][3]=	-7	;
assign conv3_kernel[2][1][4][4]=	-1	;
assign conv3_kernel[3][0][0][0]=	10	;
assign conv3_kernel[3][0][0][1]=	-16	;
assign conv3_kernel[3][0][0][2]=	13	;
assign conv3_kernel[3][0][0][3]=	-13	;
assign conv3_kernel[3][0][0][4]=	-20	;
assign conv3_kernel[3][0][1][0]=	22	;
assign conv3_kernel[3][0][1][1]=	-11	;
assign conv3_kernel[3][0][1][2]=	0	;
assign conv3_kernel[3][0][1][3]=	1	;
assign conv3_kernel[3][0][1][4]=	34	;
assign conv3_kernel[3][0][2][0]=	-1	;
assign conv3_kernel[3][0][2][1]=	-32	;
assign conv3_kernel[3][0][2][2]=	1	;
assign conv3_kernel[3][0][2][3]=	26	;
assign conv3_kernel[3][0][2][4]=	17	;
assign conv3_kernel[3][0][3][0]=	-20	;
assign conv3_kernel[3][0][3][1]=	-9	;
assign conv3_kernel[3][0][3][2]=	16	;
assign conv3_kernel[3][0][3][3]=	-58	;
assign conv3_kernel[3][0][3][4]=	-9	;
assign conv3_kernel[3][0][4][0]=	33	;
assign conv3_kernel[3][0][4][1]=	19	;
assign conv3_kernel[3][0][4][2]=	29	;
assign conv3_kernel[3][0][4][3]=	-7	;
assign conv3_kernel[3][0][4][4]=	-32	;
assign conv3_kernel[3][1][0][0]=	17	;
assign conv3_kernel[3][1][0][1]=	8	;
assign conv3_kernel[3][1][0][2]=	8	;
assign conv3_kernel[3][1][0][3]=	-40	;
assign conv3_kernel[3][1][0][4]=	17	;
assign conv3_kernel[3][1][1][0]=	-13	;
assign conv3_kernel[3][1][1][1]=	2	;
assign conv3_kernel[3][1][1][2]=	16	;
assign conv3_kernel[3][1][1][3]=	12	;
assign conv3_kernel[3][1][1][4]=	-6	;
assign conv3_kernel[3][1][2][0]=	-16	;
assign conv3_kernel[3][1][2][1]=	0	;
assign conv3_kernel[3][1][2][2]=	59	;
assign conv3_kernel[3][1][2][3]=	42	;
assign conv3_kernel[3][1][2][4]=	29	;
assign conv3_kernel[3][1][3][0]=	66	;
assign conv3_kernel[3][1][3][1]=	-8	;
assign conv3_kernel[3][1][3][2]=	-9	;
assign conv3_kernel[3][1][3][3]=	19	;
assign conv3_kernel[3][1][3][4]=	55	;
assign conv3_kernel[3][1][4][0]=	-121	;
assign conv3_kernel[3][1][4][1]=	-13	;
assign conv3_kernel[3][1][4][2]=	11	;
assign conv3_kernel[3][1][4][3]=	12	;
assign conv3_kernel[3][1][4][4]=	-12	;
assign conv3_kernel[4][0][0][0]=	-8	;
assign conv3_kernel[4][0][0][1]=	32	;
assign conv3_kernel[4][0][0][2]=	50	;
assign conv3_kernel[4][0][0][3]=	78	;
assign conv3_kernel[4][0][0][4]=	50	;
assign conv3_kernel[4][0][1][0]=	10	;
assign conv3_kernel[4][0][1][1]=	4	;
assign conv3_kernel[4][0][1][2]=	5	;
assign conv3_kernel[4][0][1][3]=	11	;
assign conv3_kernel[4][0][1][4]=	24	;
assign conv3_kernel[4][0][2][0]=	-25	;
assign conv3_kernel[4][0][2][1]=	-8	;
assign conv3_kernel[4][0][2][2]=	22	;
assign conv3_kernel[4][0][2][3]=	-36	;
assign conv3_kernel[4][0][2][4]=	-45	;
assign conv3_kernel[4][0][3][0]=	-10	;
assign conv3_kernel[4][0][3][1]=	1	;
assign conv3_kernel[4][0][3][2]=	37	;
assign conv3_kernel[4][0][3][3]=	-24	;
assign conv3_kernel[4][0][3][4]=	-1	;
assign conv3_kernel[4][0][4][0]=	9	;
assign conv3_kernel[4][0][4][1]=	-11	;
assign conv3_kernel[4][0][4][2]=	20	;
assign conv3_kernel[4][0][4][3]=	5	;
assign conv3_kernel[4][0][4][4]=	-29	;
assign conv3_kernel[4][1][0][0]=	22	;
assign conv3_kernel[4][1][0][1]=	-15	;
assign conv3_kernel[4][1][0][2]=	-34	;
assign conv3_kernel[4][1][0][3]=	-75	;
assign conv3_kernel[4][1][0][4]=	-18	;
assign conv3_kernel[4][1][1][0]=	-21	;
assign conv3_kernel[4][1][1][1]=	-13	;
assign conv3_kernel[4][1][1][2]=	-7	;
assign conv3_kernel[4][1][1][3]=	14	;
assign conv3_kernel[4][1][1][4]=	73	;
assign conv3_kernel[4][1][2][0]=	-37	;
assign conv3_kernel[4][1][2][1]=	6	;
assign conv3_kernel[4][1][2][2]=	31	;
assign conv3_kernel[4][1][2][3]=	50	;
assign conv3_kernel[4][1][2][4]=	48	;
assign conv3_kernel[4][1][3][0]=	-3	;
assign conv3_kernel[4][1][3][1]=	33	;
assign conv3_kernel[4][1][3][2]=	5	;
assign conv3_kernel[4][1][3][3]=	18	;
assign conv3_kernel[4][1][3][4]=	-10	;
assign conv3_kernel[4][1][4][0]=	-35	;
assign conv3_kernel[4][1][4][1]=	23	;
assign conv3_kernel[4][1][4][2]=	12	;
assign conv3_kernel[4][1][4][3]=	26	;
assign conv3_kernel[4][1][4][4]=	-3	;
assign conv3_kernel[5][0][0][0]=	77	;
assign conv3_kernel[5][0][0][1]=	33	;
assign conv3_kernel[5][0][0][2]=	23	;
assign conv3_kernel[5][0][0][3]=	-17	;
assign conv3_kernel[5][0][0][4]=	-34	;
assign conv3_kernel[5][0][1][0]=	45	;
assign conv3_kernel[5][0][1][1]=	12	;
assign conv3_kernel[5][0][1][2]=	4	;
assign conv3_kernel[5][0][1][3]=	-3	;
assign conv3_kernel[5][0][1][4]=	8	;
assign conv3_kernel[5][0][2][0]=	15	;
assign conv3_kernel[5][0][2][1]=	-6	;
assign conv3_kernel[5][0][2][2]=	-9	;
assign conv3_kernel[5][0][2][3]=	3	;
assign conv3_kernel[5][0][2][4]=	-22	;
assign conv3_kernel[5][0][3][0]=	0	;
assign conv3_kernel[5][0][3][1]=	13	;
assign conv3_kernel[5][0][3][2]=	-9	;
assign conv3_kernel[5][0][3][3]=	-3	;
assign conv3_kernel[5][0][3][4]=	-2	;
assign conv3_kernel[5][0][4][0]=	3	;
assign conv3_kernel[5][0][4][1]=	-23	;
assign conv3_kernel[5][0][4][2]=	-23	;
assign conv3_kernel[5][0][4][3]=	8	;
assign conv3_kernel[5][0][4][4]=	-34	;
assign conv3_kernel[5][1][0][0]=	-44	;
assign conv3_kernel[5][1][0][1]=	5	;
assign conv3_kernel[5][1][0][2]=	16	;
assign conv3_kernel[5][1][0][3]=	-3	;
assign conv3_kernel[5][1][0][4]=	6	;
assign conv3_kernel[5][1][1][0]=	-18	;
assign conv3_kernel[5][1][1][1]=	31	;
assign conv3_kernel[5][1][1][2]=	12	;
assign conv3_kernel[5][1][1][3]=	21	;
assign conv3_kernel[5][1][1][4]=	9	;
assign conv3_kernel[5][1][2][0]=	61	;
assign conv3_kernel[5][1][2][1]=	-7	;
assign conv3_kernel[5][1][2][2]=	2	;
assign conv3_kernel[5][1][2][3]=	18	;
assign conv3_kernel[5][1][2][4]=	37	;
assign conv3_kernel[5][1][3][0]=	96	;
assign conv3_kernel[5][1][3][1]=	12	;
assign conv3_kernel[5][1][3][2]=	-13	;
assign conv3_kernel[5][1][3][3]=	24	;
assign conv3_kernel[5][1][3][4]=	10	;
assign conv3_kernel[5][1][4][0]=	84	;
assign conv3_kernel[5][1][4][1]=	25	;
assign conv3_kernel[5][1][4][2]=	19	;
assign conv3_kernel[5][1][4][3]=	2	;
assign conv3_kernel[5][1][4][4]=	-21	;
assign conv3_kernel[6][0][0][0]=	-11	;
assign conv3_kernel[6][0][0][1]=	-47	;
assign conv3_kernel[6][0][0][2]=	-24	;
assign conv3_kernel[6][0][0][3]=	6	;
assign conv3_kernel[6][0][0][4]=	35	;
assign conv3_kernel[6][0][1][0]=	-15	;
assign conv3_kernel[6][0][1][1]=	17	;
assign conv3_kernel[6][0][1][2]=	9	;
assign conv3_kernel[6][0][1][3]=	9	;
assign conv3_kernel[6][0][1][4]=	23	;
assign conv3_kernel[6][0][2][0]=	17	;
assign conv3_kernel[6][0][2][1]=	-2	;
assign conv3_kernel[6][0][2][2]=	-14	;
assign conv3_kernel[6][0][2][3]=	58	;
assign conv3_kernel[6][0][2][4]=	18	;
assign conv3_kernel[6][0][3][0]=	-8	;
assign conv3_kernel[6][0][3][1]=	18	;
assign conv3_kernel[6][0][3][2]=	-6	;
assign conv3_kernel[6][0][3][3]=	24	;
assign conv3_kernel[6][0][3][4]=	38	;
assign conv3_kernel[6][0][4][0]=	30	;
assign conv3_kernel[6][0][4][1]=	-11	;
assign conv3_kernel[6][0][4][2]=	0	;
assign conv3_kernel[6][0][4][3]=	9	;
assign conv3_kernel[6][0][4][4]=	-9	;
assign conv3_kernel[6][1][0][0]=	44	;
assign conv3_kernel[6][1][0][1]=	8	;
assign conv3_kernel[6][1][0][2]=	-31	;
assign conv3_kernel[6][1][0][3]=	-72	;
assign conv3_kernel[6][1][0][4]=	-37	;
assign conv3_kernel[6][1][1][0]=	-20	;
assign conv3_kernel[6][1][1][1]=	2	;
assign conv3_kernel[6][1][1][2]=	-6	;
assign conv3_kernel[6][1][1][3]=	-11	;
assign conv3_kernel[6][1][1][4]=	-9	;
assign conv3_kernel[6][1][2][0]=	39	;
assign conv3_kernel[6][1][2][1]=	13	;
assign conv3_kernel[6][1][2][2]=	18	;
assign conv3_kernel[6][1][2][3]=	68	;
assign conv3_kernel[6][1][2][4]=	10	;
assign conv3_kernel[6][1][3][0]=	45	;
assign conv3_kernel[6][1][3][1]=	15	;
assign conv3_kernel[6][1][3][2]=	9	;
assign conv3_kernel[6][1][3][3]=	22	;
assign conv3_kernel[6][1][3][4]=	49	;
assign conv3_kernel[6][1][4][0]=	-31	;
assign conv3_kernel[6][1][4][1]=	-15	;
assign conv3_kernel[6][1][4][2]=	-11	;
assign conv3_kernel[6][1][4][3]=	-39	;
assign conv3_kernel[6][1][4][4]=	22	;
assign conv3_kernel[7][0][0][0]=	-15	;
assign conv3_kernel[7][0][0][1]=	-1	;
assign conv3_kernel[7][0][0][2]=	-41	;
assign conv3_kernel[7][0][0][3]=	-22	;
assign conv3_kernel[7][0][0][4]=	-4	;
assign conv3_kernel[7][0][1][0]=	-71	;
assign conv3_kernel[7][0][1][1]=	4	;
assign conv3_kernel[7][0][1][2]=	18	;
assign conv3_kernel[7][0][1][3]=	9	;
assign conv3_kernel[7][0][1][4]=	4	;
assign conv3_kernel[7][0][2][0]=	13	;
assign conv3_kernel[7][0][2][1]=	12	;
assign conv3_kernel[7][0][2][2]=	9	;
assign conv3_kernel[7][0][2][3]=	7	;
assign conv3_kernel[7][0][2][4]=	16	;
assign conv3_kernel[7][0][3][0]=	25	;
assign conv3_kernel[7][0][3][1]=	3	;
assign conv3_kernel[7][0][3][2]=	-2	;
assign conv3_kernel[7][0][3][3]=	-23	;
assign conv3_kernel[7][0][3][4]=	-62	;
assign conv3_kernel[7][0][4][0]=	-2	;
assign conv3_kernel[7][0][4][1]=	2	;
assign conv3_kernel[7][0][4][2]=	-14	;
assign conv3_kernel[7][0][4][3]=	6	;
assign conv3_kernel[7][0][4][4]=	33	;
assign conv3_kernel[7][1][0][0]=	10	;
assign conv3_kernel[7][1][0][1]=	40	;
assign conv3_kernel[7][1][0][2]=	5	;
assign conv3_kernel[7][1][0][3]=	2	;
assign conv3_kernel[7][1][0][4]=	35	;
assign conv3_kernel[7][1][1][0]=	39	;
assign conv3_kernel[7][1][1][1]=	5	;
assign conv3_kernel[7][1][1][2]=	8	;
assign conv3_kernel[7][1][1][3]=	9	;
assign conv3_kernel[7][1][1][4]=	15	;
assign conv3_kernel[7][1][2][0]=	-37	;
assign conv3_kernel[7][1][2][1]=	-27	;
assign conv3_kernel[7][1][2][2]=	34	;
assign conv3_kernel[7][1][2][3]=	56	;
assign conv3_kernel[7][1][2][4]=	-6	;
assign conv3_kernel[7][1][3][0]=	-23	;
assign conv3_kernel[7][1][3][1]=	24	;
assign conv3_kernel[7][1][3][2]=	35	;
assign conv3_kernel[7][1][3][3]=	21	;
assign conv3_kernel[7][1][3][4]=	-42	;
assign conv3_kernel[7][1][4][0]=	37	;
assign conv3_kernel[7][1][4][1]=	20	;
assign conv3_kernel[7][1][4][2]=	27	;
assign conv3_kernel[7][1][4][3]=	-10	;
assign conv3_kernel[7][1][4][4]=	-70	;
assign conv3_kernel[8][0][0][0]=	-76	;
assign conv3_kernel[8][0][0][1]=	-29	;
assign conv3_kernel[8][0][0][2]=	15	;
assign conv3_kernel[8][0][0][3]=	-3	;
assign conv3_kernel[8][0][0][4]=	22	;
assign conv3_kernel[8][0][1][0]=	-116	;
assign conv3_kernel[8][0][1][1]=	2	;
assign conv3_kernel[8][0][1][2]=	2	;
assign conv3_kernel[8][0][1][3]=	5	;
assign conv3_kernel[8][0][1][4]=	-8	;
assign conv3_kernel[8][0][2][0]=	22	;
assign conv3_kernel[8][0][2][1]=	-18	;
assign conv3_kernel[8][0][2][2]=	16	;
assign conv3_kernel[8][0][2][3]=	13	;
assign conv3_kernel[8][0][2][4]=	40	;
assign conv3_kernel[8][0][3][0]=	-2	;
assign conv3_kernel[8][0][3][1]=	-3	;
assign conv3_kernel[8][0][3][2]=	10	;
assign conv3_kernel[8][0][3][3]=	-15	;
assign conv3_kernel[8][0][3][4]=	-3	;
assign conv3_kernel[8][0][4][0]=	18	;
assign conv3_kernel[8][0][4][1]=	7	;
assign conv3_kernel[8][0][4][2]=	-2	;
assign conv3_kernel[8][0][4][3]=	8	;
assign conv3_kernel[8][0][4][4]=	-5	;
assign conv3_kernel[8][1][0][0]=	57	;
assign conv3_kernel[8][1][0][1]=	40	;
assign conv3_kernel[8][1][0][2]=	3	;
assign conv3_kernel[8][1][0][3]=	-6	;
assign conv3_kernel[8][1][0][4]=	30	;
assign conv3_kernel[8][1][1][0]=	25	;
assign conv3_kernel[8][1][1][1]=	7	;
assign conv3_kernel[8][1][1][2]=	10	;
assign conv3_kernel[8][1][1][3]=	27	;
assign conv3_kernel[8][1][1][4]=	31	;
assign conv3_kernel[8][1][2][0]=	6	;
assign conv3_kernel[8][1][2][1]=	-33	;
assign conv3_kernel[8][1][2][2]=	-40	;
assign conv3_kernel[8][1][2][3]=	-16	;
assign conv3_kernel[8][1][2][4]=	-32	;
assign conv3_kernel[8][1][3][0]=	-17	;
assign conv3_kernel[8][1][3][1]=	-14	;
assign conv3_kernel[8][1][3][2]=	-16	;
assign conv3_kernel[8][1][3][3]=	0	;
assign conv3_kernel[8][1][3][4]=	-27	;
assign conv3_kernel[8][1][4][0]=	-76	;
assign conv3_kernel[8][1][4][1]=	9	;
assign conv3_kernel[8][1][4][2]=	9	;
assign conv3_kernel[8][1][4][3]=	11	;
assign conv3_kernel[8][1][4][4]=	-60	;
assign conv3_kernel[9][0][0][0]=	43	;
assign conv3_kernel[9][0][0][1]=	-28	;
assign conv3_kernel[9][0][0][2]=	-28	;
assign conv3_kernel[9][0][0][3]=	-49	;
assign conv3_kernel[9][0][0][4]=	-24	;
assign conv3_kernel[9][0][1][0]=	41	;
assign conv3_kernel[9][0][1][1]=	-18	;
assign conv3_kernel[9][0][1][2]=	17	;
assign conv3_kernel[9][0][1][3]=	18	;
assign conv3_kernel[9][0][1][4]=	9	;
assign conv3_kernel[9][0][2][0]=	-3	;
assign conv3_kernel[9][0][2][1]=	-14	;
assign conv3_kernel[9][0][2][2]=	70	;
assign conv3_kernel[9][0][2][3]=	41	;
assign conv3_kernel[9][0][2][4]=	0	;
assign conv3_kernel[9][0][3][0]=	-19	;
assign conv3_kernel[9][0][3][1]=	-16	;
assign conv3_kernel[9][0][3][2]=	42	;
assign conv3_kernel[9][0][3][3]=	-30	;
assign conv3_kernel[9][0][3][4]=	1	;
assign conv3_kernel[9][0][4][0]=	4	;
assign conv3_kernel[9][0][4][1]=	-38	;
assign conv3_kernel[9][0][4][2]=	44	;
assign conv3_kernel[9][0][4][3]=	24	;
assign conv3_kernel[9][0][4][4]=	-22	;
assign conv3_kernel[9][1][0][0]=	-7	;
assign conv3_kernel[9][1][0][1]=	13	;
assign conv3_kernel[9][1][0][2]=	44	;
assign conv3_kernel[9][1][0][3]=	-36	;
assign conv3_kernel[9][1][0][4]=	-8	;
assign conv3_kernel[9][1][1][0]=	-5	;
assign conv3_kernel[9][1][1][1]=	-12	;
assign conv3_kernel[9][1][1][2]=	11	;
assign conv3_kernel[9][1][1][3]=	-25	;
assign conv3_kernel[9][1][1][4]=	-35	;
assign conv3_kernel[9][1][2][0]=	-2	;
assign conv3_kernel[9][1][2][1]=	-12	;
assign conv3_kernel[9][1][2][2]=	29	;
assign conv3_kernel[9][1][2][3]=	-3	;
assign conv3_kernel[9][1][2][4]=	-1	;
assign conv3_kernel[9][1][3][0]=	17	;
assign conv3_kernel[9][1][3][1]=	7	;
assign conv3_kernel[9][1][3][2]=	4	;
assign conv3_kernel[9][1][3][3]=	4	;
assign conv3_kernel[9][1][3][4]=	3	;
assign conv3_kernel[9][1][4][0]=	14	;
assign conv3_kernel[9][1][4][1]=	27	;
assign conv3_kernel[9][1][4][2]=	1	;
assign conv3_kernel[9][1][4][3]=	-4	;
assign conv3_kernel[9][1][4][4]=	-13	;
assign connect_matrix [0][0]=	-43	;
assign connect_matrix [0][1]=	49	;
assign connect_matrix [0][2]=	-7	;
assign connect_matrix [0][3]=	-39	;
assign connect_matrix [0][4]=	7	;
assign connect_matrix [0][5]=	-8	;
assign connect_matrix [0][6]=	-3	;
assign connect_matrix [0][7]=	-2	;
assign connect_matrix [0][8]=	25	;
assign connect_matrix [0][9]=	-24	;
assign connect_matrix [1][0]=	54	;
assign connect_matrix [1][1]=	-18	;
assign connect_matrix [1][2]=	-51	;
assign connect_matrix [1][3]=	-39	;
assign connect_matrix [1][4]=	0	;
assign connect_matrix [1][5]=	19	;
assign connect_matrix [1][6]=	20	;
assign connect_matrix [1][7]=	-94	;
assign connect_matrix [1][8]=	50	;
assign connect_matrix [1][9]=	74	;
assign connect_matrix [2][0]=	20	;
assign connect_matrix [2][1]=	42	;
assign connect_matrix [2][2]=	-2	;
assign connect_matrix [2][3]=	19	;
assign connect_matrix [2][4]=	-45	;
assign connect_matrix [2][5]=	24	;
assign connect_matrix [2][6]=	6	;
assign connect_matrix [2][7]=	-22	;
assign connect_matrix [2][8]=	-57	;
assign connect_matrix [2][9]=	-3	;
assign connect_matrix [3][0]=	-14	;
assign connect_matrix [3][1]=	-2	;
assign connect_matrix [3][2]=	-32	;
assign connect_matrix [3][3]=	-1	;
assign connect_matrix [3][4]=	-9	;
assign connect_matrix [3][5]=	47	;
assign connect_matrix [3][6]=	-13	;
assign connect_matrix [3][7]=	22	;
assign connect_matrix [3][8]=	-45	;
assign connect_matrix [3][9]=	22	;
assign connect_matrix [4][0]=	0	;
assign connect_matrix [4][1]=	-18	;
assign connect_matrix [4][2]=	-5	;
assign connect_matrix [4][3]=	-17	;
assign connect_matrix [4][4]=	-34	;
assign connect_matrix [4][5]=	-46	;
assign connect_matrix [4][6]=	64	;
assign connect_matrix [4][7]=	28	;
assign connect_matrix [4][8]=	-20	;
assign connect_matrix [4][9]=	23	;
assign connect_matrix [5][0]=	18	;
assign connect_matrix [5][1]=	-32	;
assign connect_matrix [5][2]=	-34	;
assign connect_matrix [5][3]=	-13	;
assign connect_matrix [5][4]=	42	;
assign connect_matrix [5][5]=	25	;
assign connect_matrix [5][6]=	-7	;
assign connect_matrix [5][7]=	20	;
assign connect_matrix [5][8]=	-6	;
assign connect_matrix [5][9]=	-38	;
assign connect_matrix [6][0]=	-52	;
assign connect_matrix [6][1]=	26	;
assign connect_matrix [6][2]=	21	;
assign connect_matrix [6][3]=	9	;
assign connect_matrix [6][4]=	62	;
assign connect_matrix [6][5]=	-91	;
assign connect_matrix [6][6]=	13	;
assign connect_matrix [6][7]=	-14	;
assign connect_matrix [6][8]=	-14	;
assign connect_matrix [6][9]=	-16	;
assign connect_matrix [7][0]=	-32	;
assign connect_matrix [7][1]=	-43	;
assign connect_matrix [7][2]=	54	;
assign connect_matrix [7][3]=	20	;
assign connect_matrix [7][4]=	-5	;
assign connect_matrix [7][5]=	28	;
assign connect_matrix [7][6]=	0	;
assign connect_matrix [7][7]=	-39	;
assign connect_matrix [7][8]=	27	;
assign connect_matrix [7][9]=	17	;
assign connect_matrix [8][0]=	7	;
assign connect_matrix [8][1]=	-2	;
assign connect_matrix [8][2]=	2	;
assign connect_matrix [8][3]=	58	;
assign connect_matrix [8][4]=	-14	;
assign connect_matrix [8][5]=	-9	;
assign connect_matrix [8][6]=	-29	;
assign connect_matrix [8][7]=	12	;
assign connect_matrix [8][8]=	11	;
assign connect_matrix [8][9]=	-9	;
assign connect_matrix [9][0]=	27	;
assign connect_matrix [9][1]=	-7	;
assign connect_matrix [9][2]=	38	;
assign connect_matrix [9][3]=	-20	;
assign connect_matrix [9][4]=	-11	;
assign connect_matrix [9][5]=	-23	;
assign connect_matrix [9][6]=	-35	;
assign connect_matrix [9][7]=	42	;
assign connect_matrix [9][8]=	-31	;
assign connect_matrix [9][9]=	17	;






// end
//     end
// endmodule