// module kernel_matrix_trained(conv1_kernel,conv2_kernel,conv3_kernel,connect_matrix);
//     parameter bitwidth=32;
//     output reg signed [bitwidth-1:0] conv1_kernel [1:0][4:0][4:0];
// 	output reg signed [bitwidth-1:0] conv2_kernel [1:0][1:0][4:0][4:0];
// 	output reg signed [bitwidth-1:0] conv3_kernel [9:0][1:0][4:0][4:0];
// 	output reg signed [bitwidth-1:0] connect_matrix [9:0][9:0];
//     always@(*) begin
initial begin
conv1_kernel[0][0][0]=	-37426	;
conv1_kernel[0][0][1]=	-25898	;
conv1_kernel[0][0][2]=	11740	;
conv1_kernel[0][0][3]=	-6400	;
conv1_kernel[0][0][4]=	13650	;
conv1_kernel[0][1][0]=	-45961	;
conv1_kernel[0][1][1]=	12264	;
conv1_kernel[0][1][2]=	11523	;
conv1_kernel[0][1][3]=	11971	;
conv1_kernel[0][1][4]=	6510	;
conv1_kernel[0][2][0]=	-36322	;
conv1_kernel[0][2][1]=	35186	;
conv1_kernel[0][2][2]=	19545	;
conv1_kernel[0][2][3]=	18770	;
conv1_kernel[0][2][4]=	-2499	;
conv1_kernel[0][3][0]=	-13884	;
conv1_kernel[0][3][1]=	7890	;
conv1_kernel[0][3][2]=	16199	;
conv1_kernel[0][3][3]=	8499	;
conv1_kernel[0][3][4]=	2267	;
conv1_kernel[0][4][0]=	-9035	;
conv1_kernel[0][4][1]=	17393	;
conv1_kernel[0][4][2]=	-3303	;
conv1_kernel[0][4][3]=	-7284	;
conv1_kernel[0][4][4]=	-18060	;
conv1_kernel[1][0][0]=	7158	;
conv1_kernel[1][0][1]=	2280	;
conv1_kernel[1][0][2]=	3476	;
conv1_kernel[1][0][3]=	-6045	;
conv1_kernel[1][0][4]=	-8221	;
conv1_kernel[1][1][0]=	13526	;
conv1_kernel[1][1][1]=	4535	;
conv1_kernel[1][1][2]=	-975	;
conv1_kernel[1][1][3]=	277	;
conv1_kernel[1][1][4]=	-1929	;
conv1_kernel[1][2][0]=	11894	;
conv1_kernel[1][2][1]=	14499	;
conv1_kernel[1][2][2]=	1099	;
conv1_kernel[1][2][3]=	242	;
conv1_kernel[1][2][4]=	15540	;
conv1_kernel[1][3][0]=	-3193	;
conv1_kernel[1][3][1]=	21456	;
conv1_kernel[1][3][2]=	34254	;
conv1_kernel[1][3][3]=	14447	;
conv1_kernel[1][3][4]=	3232	;
conv1_kernel[1][4][0]=	-130	;
conv1_kernel[1][4][1]=	-2939	;
conv1_kernel[1][4][2]=	1024	;
conv1_kernel[1][4][3]=	7644	;
conv1_kernel[1][4][4]=	7933	;
conv2_kernel[0][0][0][0]=	11357	;
conv2_kernel[0][0][0][1]=	27553	;
conv2_kernel[0][0][0][2]=	35193	;
conv2_kernel[0][0][0][3]=	-110	;
conv2_kernel[0][0][0][4]=	-3063	;
conv2_kernel[0][0][1][0]=	-35933	;
conv2_kernel[0][0][1][1]=	25526	;
conv2_kernel[0][0][1][2]=	17952	;
conv2_kernel[0][0][1][3]=	-11616	;
conv2_kernel[0][0][1][4]=	-12050	;
conv2_kernel[0][0][2][0]=	8202	;
conv2_kernel[0][0][2][1]=	-14823	;
conv2_kernel[0][0][2][2]=	-5051	;
conv2_kernel[0][0][2][3]=	3265	;
conv2_kernel[0][0][2][4]=	22981	;
conv2_kernel[0][0][3][0]=	14209	;
conv2_kernel[0][0][3][1]=	2477	;
conv2_kernel[0][0][3][2]=	-570	;
conv2_kernel[0][0][3][3]=	30513	;
conv2_kernel[0][0][3][4]=	11196	;
conv2_kernel[0][0][4][0]=	1273	;
conv2_kernel[0][0][4][1]=	-30923	;
conv2_kernel[0][0][4][2]=	-40251	;
conv2_kernel[0][0][4][3]=	-58296	;
conv2_kernel[0][0][4][4]=	-8594	;
conv2_kernel[0][1][0][0]=	-31034	;
conv2_kernel[0][1][0][1]=	-14823	;
conv2_kernel[0][1][0][2]=	4066	;
conv2_kernel[0][1][0][3]=	16529	;
conv2_kernel[0][1][0][4]=	-28052	;
conv2_kernel[0][1][1][0]=	-41733	;
conv2_kernel[0][1][1][1]=	27	;
conv2_kernel[0][1][1][2]=	3188	;
conv2_kernel[0][1][1][3]=	13532	;
conv2_kernel[0][1][1][4]=	31654	;
conv2_kernel[0][1][2][0]=	32339	;
conv2_kernel[0][1][2][1]=	59865	;
conv2_kernel[0][1][2][2]=	70248	;
conv2_kernel[0][1][2][3]=	81100	;
conv2_kernel[0][1][2][4]=	23545	;
conv2_kernel[0][1][3][0]=	-18207	;
conv2_kernel[0][1][3][1]=	-27417	;
conv2_kernel[0][1][3][2]=	-747	;
conv2_kernel[0][1][3][3]=	-30673	;
conv2_kernel[0][1][3][4]=	-92763	;
conv2_kernel[0][1][4][0]=	-8852	;
conv2_kernel[0][1][4][1]=	9747	;
conv2_kernel[0][1][4][2]=	-29886	;
conv2_kernel[0][1][4][3]=	-46309	;
conv2_kernel[0][1][4][4]=	1451	;
conv2_kernel[1][0][0][0]=	41474	;
conv2_kernel[1][0][0][1]=	28551	;
conv2_kernel[1][0][0][2]=	-15185	;
conv2_kernel[1][0][0][3]=	-30910	;
conv2_kernel[1][0][0][4]=	-12179	;
conv2_kernel[1][0][1][0]=	-34642	;
conv2_kernel[1][0][1][1]=	-47993	;
conv2_kernel[1][0][1][2]=	28240	;
conv2_kernel[1][0][1][3]=	-2252	;
conv2_kernel[1][0][1][4]=	-29528	;
conv2_kernel[1][0][2][0]=	-38238	;
conv2_kernel[1][0][2][1]=	-34596	;
conv2_kernel[1][0][2][2]=	23584	;
conv2_kernel[1][0][2][3]=	25081	;
conv2_kernel[1][0][2][4]=	11846	;
conv2_kernel[1][0][3][0]=	9781	;
conv2_kernel[1][0][3][1]=	-20544	;
conv2_kernel[1][0][3][2]=	-63142	;
conv2_kernel[1][0][3][3]=	-3533	;
conv2_kernel[1][0][3][4]=	4149	;
conv2_kernel[1][0][4][0]=	15554	;
conv2_kernel[1][0][4][1]=	8455	;
conv2_kernel[1][0][4][2]=	6250	;
conv2_kernel[1][0][4][3]=	-2677	;
conv2_kernel[1][0][4][4]=	3772	;
conv2_kernel[1][1][0][0]=	-48717	;
conv2_kernel[1][1][0][1]=	-33008	;
conv2_kernel[1][1][0][2]=	-42483	;
conv2_kernel[1][1][0][3]=	-43827	;
conv2_kernel[1][1][0][4]=	-49536	;
conv2_kernel[1][1][1][0]=	-11933	;
conv2_kernel[1][1][1][1]=	-60122	;
conv2_kernel[1][1][1][2]=	10607	;
conv2_kernel[1][1][1][3]=	19349	;
conv2_kernel[1][1][1][4]=	36363	;
conv2_kernel[1][1][2][0]=	127225	;
conv2_kernel[1][1][2][1]=	110339	;
conv2_kernel[1][1][2][2]=	48267	;
conv2_kernel[1][1][2][3]=	4906	;
conv2_kernel[1][1][2][4]=	35826	;
conv2_kernel[1][1][3][0]=	-50913	;
conv2_kernel[1][1][3][1]=	16707	;
conv2_kernel[1][1][3][2]=	124	;
conv2_kernel[1][1][3][3]=	15023	;
conv2_kernel[1][1][3][4]=	-11326	;
conv2_kernel[1][1][4][0]=	-74539	;
conv2_kernel[1][1][4][1]=	-13160	;
conv2_kernel[1][1][4][2]=	14323	;
conv2_kernel[1][1][4][3]=	10338	;
conv2_kernel[1][1][4][4]=	-3452	;
conv3_kernel[0][0][0][0]=	-66980	;
conv3_kernel[0][0][0][1]=	-15322	;
conv3_kernel[0][0][0][2]=	19481	;
conv3_kernel[0][0][0][3]=	25043	;
conv3_kernel[0][0][0][4]=	5624	;
conv3_kernel[0][0][1][0]=	-29712	;
conv3_kernel[0][0][1][1]=	-3193	;
conv3_kernel[0][0][1][2]=	5066	;
conv3_kernel[0][0][1][3]=	-6730	;
conv3_kernel[0][0][1][4]=	17886	;
conv3_kernel[0][0][2][0]=	28450	;
conv3_kernel[0][0][2][1]=	17726	;
conv3_kernel[0][0][2][2]=	20303	;
conv3_kernel[0][0][2][3]=	7414	;
conv3_kernel[0][0][2][4]=	1164	;
conv3_kernel[0][0][3][0]=	12601	;
conv3_kernel[0][0][3][1]=	-4678	;
conv3_kernel[0][0][3][2]=	32335	;
conv3_kernel[0][0][3][3]=	-23053	;
conv3_kernel[0][0][3][4]=	13738	;
conv3_kernel[0][0][4][0]=	6643	;
conv3_kernel[0][0][4][1]=	-16523	;
conv3_kernel[0][0][4][2]=	7355	;
conv3_kernel[0][0][4][3]=	1847	;
conv3_kernel[0][0][4][4]=	1316	;
conv3_kernel[0][1][0][0]=	-19694	;
conv3_kernel[0][1][0][1]=	20404	;
conv3_kernel[0][1][0][2]=	14137	;
conv3_kernel[0][1][0][3]=	-36355	;
conv3_kernel[0][1][0][4]=	-17801	;
conv3_kernel[0][1][1][0]=	-73557	;
conv3_kernel[0][1][1][1]=	5970	;
conv3_kernel[0][1][1][2]=	22645	;
conv3_kernel[0][1][1][3]=	2247	;
conv3_kernel[0][1][1][4]=	-2265	;
conv3_kernel[0][1][2][0]=	-49179	;
conv3_kernel[0][1][2][1]=	-4379	;
conv3_kernel[0][1][2][2]=	27997	;
conv3_kernel[0][1][2][3]=	25622	;
conv3_kernel[0][1][2][4]=	-48223	;
conv3_kernel[0][1][3][0]=	54548	;
conv3_kernel[0][1][3][1]=	3118	;
conv3_kernel[0][1][3][2]=	-3068	;
conv3_kernel[0][1][3][3]=	-17141	;
conv3_kernel[0][1][3][4]=	25193	;
conv3_kernel[0][1][4][0]=	84191	;
conv3_kernel[0][1][4][1]=	-20419	;
conv3_kernel[0][1][4][2]=	3787	;
conv3_kernel[0][1][4][3]=	13358	;
conv3_kernel[0][1][4][4]=	51081	;
conv3_kernel[1][0][0][0]=	37917	;
conv3_kernel[1][0][0][1]=	19369	;
conv3_kernel[1][0][0][2]=	-5439	;
conv3_kernel[1][0][0][3]=	-14253	;
conv3_kernel[1][0][0][4]=	-84718	;
conv3_kernel[1][0][1][0]=	12729	;
conv3_kernel[1][0][1][1]=	12323	;
conv3_kernel[1][0][1][2]=	-11850	;
conv3_kernel[1][0][1][3]=	-3913	;
conv3_kernel[1][0][1][4]=	-82811	;
conv3_kernel[1][0][2][0]=	-51385	;
conv3_kernel[1][0][2][1]=	-11353	;
conv3_kernel[1][0][2][2]=	-698	;
conv3_kernel[1][0][2][3]=	2501	;
conv3_kernel[1][0][2][4]=	54857	;
conv3_kernel[1][0][3][0]=	-25352	;
conv3_kernel[1][0][3][1]=	29117	;
conv3_kernel[1][0][3][2]=	40040	;
conv3_kernel[1][0][3][3]=	-1051	;
conv3_kernel[1][0][3][4]=	42370	;
conv3_kernel[1][0][4][0]=	40154	;
conv3_kernel[1][0][4][1]=	38235	;
conv3_kernel[1][0][4][2]=	-8335	;
conv3_kernel[1][0][4][3]=	-10800	;
conv3_kernel[1][0][4][4]=	-4983	;
conv3_kernel[1][1][0][0]=	-26503	;
conv3_kernel[1][1][0][1]=	-25511	;
conv3_kernel[1][1][0][2]=	-11894	;
conv3_kernel[1][1][0][3]=	-6742	;
conv3_kernel[1][1][0][4]=	23481	;
conv3_kernel[1][1][1][0]=	21690	;
conv3_kernel[1][1][1][1]=	-5991	;
conv3_kernel[1][1][1][2]=	-20393	;
conv3_kernel[1][1][1][3]=	24611	;
conv3_kernel[1][1][1][4]=	13796	;
conv3_kernel[1][1][2][0]=	25848	;
conv3_kernel[1][1][2][1]=	7232	;
conv3_kernel[1][1][2][2]=	-14620	;
conv3_kernel[1][1][2][3]=	35113	;
conv3_kernel[1][1][2][4]=	-16831	;
conv3_kernel[1][1][3][0]=	-35753	;
conv3_kernel[1][1][3][1]=	26829	;
conv3_kernel[1][1][3][2]=	-12722	;
conv3_kernel[1][1][3][3]=	-5669	;
conv3_kernel[1][1][3][4]=	16852	;
conv3_kernel[1][1][4][0]=	-91898	;
conv3_kernel[1][1][4][1]=	21338	;
conv3_kernel[1][1][4][2]=	14528	;
conv3_kernel[1][1][4][3]=	44465	;
conv3_kernel[1][1][4][4]=	40433	;
conv3_kernel[2][0][0][0]=	30645	;
conv3_kernel[2][0][0][1]=	42773	;
conv3_kernel[2][0][0][2]=	-16359	;
conv3_kernel[2][0][0][3]=	17930	;
conv3_kernel[2][0][0][4]=	-37702	;
conv3_kernel[2][0][1][0]=	-16133	;
conv3_kernel[2][0][1][1]=	14252	;
conv3_kernel[2][0][1][2]=	9836	;
conv3_kernel[2][0][1][3]=	-2902	;
conv3_kernel[2][0][1][4]=	-44248	;
conv3_kernel[2][0][2][0]=	7610	;
conv3_kernel[2][0][2][1]=	7658	;
conv3_kernel[2][0][2][2]=	-11494	;
conv3_kernel[2][0][2][3]=	60507	;
conv3_kernel[2][0][2][4]=	35542	;
conv3_kernel[2][0][3][0]=	9282	;
conv3_kernel[2][0][3][1]=	-1949	;
conv3_kernel[2][0][3][2]=	2013	;
conv3_kernel[2][0][3][3]=	60301	;
conv3_kernel[2][0][3][4]=	17844	;
conv3_kernel[2][0][4][0]=	-6595	;
conv3_kernel[2][0][4][1]=	-22025	;
conv3_kernel[2][0][4][2]=	-30613	;
conv3_kernel[2][0][4][3]=	-3777	;
conv3_kernel[2][0][4][4]=	15325	;
conv3_kernel[2][1][0][0]=	-1587	;
conv3_kernel[2][1][0][1]=	92	;
conv3_kernel[2][1][0][2]=	8022	;
conv3_kernel[2][1][0][3]=	-260	;
conv3_kernel[2][1][0][4]=	15211	;
conv3_kernel[2][1][1][0]=	29510	;
conv3_kernel[2][1][1][1]=	10332	;
conv3_kernel[2][1][1][2]=	11439	;
conv3_kernel[2][1][1][3]=	29534	;
conv3_kernel[2][1][1][4]=	9864	;
conv3_kernel[2][1][2][0]=	-25028	;
conv3_kernel[2][1][2][1]=	-6160	;
conv3_kernel[2][1][2][2]=	9530	;
conv3_kernel[2][1][2][3]=	48239	;
conv3_kernel[2][1][2][4]=	-45946	;
conv3_kernel[2][1][3][0]=	-7204	;
conv3_kernel[2][1][3][1]=	6793	;
conv3_kernel[2][1][3][2]=	15615	;
conv3_kernel[2][1][3][3]=	-30731	;
conv3_kernel[2][1][3][4]=	-35546	;
conv3_kernel[2][1][4][0]=	25684	;
conv3_kernel[2][1][4][1]=	-16287	;
conv3_kernel[2][1][4][2]=	-34701	;
conv3_kernel[2][1][4][3]=	-6919	;
conv3_kernel[2][1][4][4]=	-1217	;
conv3_kernel[3][0][0][0]=	10291	;
conv3_kernel[3][0][0][1]=	-16341	;
conv3_kernel[3][0][0][2]=	12996	;
conv3_kernel[3][0][0][3]=	-13710	;
conv3_kernel[3][0][0][4]=	-20665	;
conv3_kernel[3][0][1][0]=	22260	;
conv3_kernel[3][0][1][1]=	-11472	;
conv3_kernel[3][0][1][2]=	-470	;
conv3_kernel[3][0][1][3]=	1214	;
conv3_kernel[3][0][1][4]=	35253	;
conv3_kernel[3][0][2][0]=	-747	;
conv3_kernel[3][0][2][1]=	-32622	;
conv3_kernel[3][0][2][2]=	574	;
conv3_kernel[3][0][2][3]=	26201	;
conv3_kernel[3][0][2][4]=	17754	;
conv3_kernel[3][0][3][0]=	-20013	;
conv3_kernel[3][0][3][1]=	-9373	;
conv3_kernel[3][0][3][2]=	16870	;
conv3_kernel[3][0][3][3]=	-59902	;
conv3_kernel[3][0][3][4]=	-9479	;
conv3_kernel[3][0][4][0]=	33529	;
conv3_kernel[3][0][4][1]=	19839	;
conv3_kernel[3][0][4][2]=	30047	;
conv3_kernel[3][0][4][3]=	-6782	;
conv3_kernel[3][0][4][4]=	-32650	;
conv3_kernel[3][1][0][0]=	17059	;
conv3_kernel[3][1][0][1]=	8232	;
conv3_kernel[3][1][0][2]=	8535	;
conv3_kernel[3][1][0][3]=	-41227	;
conv3_kernel[3][1][0][4]=	17573	;
conv3_kernel[3][1][1][0]=	-13430	;
conv3_kernel[3][1][1][1]=	1852	;
conv3_kernel[3][1][1][2]=	16118	;
conv3_kernel[3][1][1][3]=	12704	;
conv3_kernel[3][1][1][4]=	-6624	;
conv3_kernel[3][1][2][0]=	-16189	;
conv3_kernel[3][1][2][1]=	67	;
conv3_kernel[3][1][2][2]=	60734	;
conv3_kernel[3][1][2][3]=	43357	;
conv3_kernel[3][1][2][4]=	29893	;
conv3_kernel[3][1][3][0]=	67453	;
conv3_kernel[3][1][3][1]=	-8259	;
conv3_kernel[3][1][3][2]=	-9518	;
conv3_kernel[3][1][3][3]=	19306	;
conv3_kernel[3][1][3][4]=	55900	;
conv3_kernel[3][1][4][0]=	-123942	;
conv3_kernel[3][1][4][1]=	-13497	;
conv3_kernel[3][1][4][2]=	11714	;
conv3_kernel[3][1][4][3]=	12740	;
conv3_kernel[3][1][4][4]=	-11780	;
conv3_kernel[4][0][0][0]=	-7791	;
conv3_kernel[4][0][0][1]=	32962	;
conv3_kernel[4][0][0][2]=	50726	;
conv3_kernel[4][0][0][3]=	79733	;
conv3_kernel[4][0][0][4]=	50857	;
conv3_kernel[4][0][1][0]=	9757	;
conv3_kernel[4][0][1][1]=	3783	;
conv3_kernel[4][0][1][2]=	5589	;
conv3_kernel[4][0][1][3]=	11516	;
conv3_kernel[4][0][1][4]=	24700	;
conv3_kernel[4][0][2][0]=	-25817	;
conv3_kernel[4][0][2][1]=	-7822	;
conv3_kernel[4][0][2][2]=	22731	;
conv3_kernel[4][0][2][3]=	-36465	;
conv3_kernel[4][0][2][4]=	-46254	;
conv3_kernel[4][0][3][0]=	-9850	;
conv3_kernel[4][0][3][1]=	1448	;
conv3_kernel[4][0][3][2]=	37616	;
conv3_kernel[4][0][3][3]=	-24316	;
conv3_kernel[4][0][3][4]=	-1091	;
conv3_kernel[4][0][4][0]=	8748	;
conv3_kernel[4][0][4][1]=	-11408	;
conv3_kernel[4][0][4][2]=	20152	;
conv3_kernel[4][0][4][3]=	5624	;
conv3_kernel[4][0][4][4]=	-29472	;
conv3_kernel[4][1][0][0]=	22095	;
conv3_kernel[4][1][0][1]=	-15612	;
conv3_kernel[4][1][0][2]=	-35054	;
conv3_kernel[4][1][0][3]=	-76876	;
conv3_kernel[4][1][0][4]=	-17920	;
conv3_kernel[4][1][1][0]=	-21556	;
conv3_kernel[4][1][1][1]=	-13733	;
conv3_kernel[4][1][1][2]=	-6823	;
conv3_kernel[4][1][1][3]=	14319	;
conv3_kernel[4][1][1][4]=	74630	;
conv3_kernel[4][1][2][0]=	-37979	;
conv3_kernel[4][1][2][1]=	6017	;
conv3_kernel[4][1][2][2]=	31395	;
conv3_kernel[4][1][2][3]=	51329	;
conv3_kernel[4][1][2][4]=	49176	;
conv3_kernel[4][1][3][0]=	-3565	;
conv3_kernel[4][1][3][1]=	33815	;
conv3_kernel[4][1][3][2]=	4857	;
conv3_kernel[4][1][3][3]=	17931	;
conv3_kernel[4][1][3][4]=	-10036	;
conv3_kernel[4][1][4][0]=	-35349	;
conv3_kernel[4][1][4][1]=	23458	;
conv3_kernel[4][1][4][2]=	12568	;
conv3_kernel[4][1][4][3]=	26252	;
conv3_kernel[4][1][4][4]=	-2683	;
conv3_kernel[5][0][0][0]=	79003	;
conv3_kernel[5][0][0][1]=	34132	;
conv3_kernel[5][0][0][2]=	23621	;
conv3_kernel[5][0][0][3]=	-17481	;
conv3_kernel[5][0][0][4]=	-34451	;
conv3_kernel[5][0][1][0]=	45580	;
conv3_kernel[5][0][1][1]=	11912	;
conv3_kernel[5][0][1][2]=	3729	;
conv3_kernel[5][0][1][3]=	-3423	;
conv3_kernel[5][0][1][4]=	8503	;
conv3_kernel[5][0][2][0]=	15192	;
conv3_kernel[5][0][2][1]=	-6307	;
conv3_kernel[5][0][2][2]=	-8984	;
conv3_kernel[5][0][2][3]=	2604	;
conv3_kernel[5][0][2][4]=	-22861	;
conv3_kernel[5][0][3][0]=	-21	;
conv3_kernel[5][0][3][1]=	13250	;
conv3_kernel[5][0][3][2]=	-9407	;
conv3_kernel[5][0][3][3]=	-2933	;
conv3_kernel[5][0][3][4]=	-2006	;
conv3_kernel[5][0][4][0]=	3280	;
conv3_kernel[5][0][4][1]=	-23992	;
conv3_kernel[5][0][4][2]=	-23538	;
conv3_kernel[5][0][4][3]=	8592	;
conv3_kernel[5][0][4][4]=	-35303	;
conv3_kernel[5][1][0][0]=	-44823	;
conv3_kernel[5][1][0][1]=	5216	;
conv3_kernel[5][1][0][2]=	16500	;
conv3_kernel[5][1][0][3]=	-2896	;
conv3_kernel[5][1][0][4]=	6030	;
conv3_kernel[5][1][1][0]=	-18283	;
conv3_kernel[5][1][1][1]=	31474	;
conv3_kernel[5][1][1][2]=	11829	;
conv3_kernel[5][1][1][3]=	21119	;
conv3_kernel[5][1][1][4]=	9160	;
conv3_kernel[5][1][2][0]=	62009	;
conv3_kernel[5][1][2][1]=	-7275	;
conv3_kernel[5][1][2][2]=	1592	;
conv3_kernel[5][1][2][3]=	18807	;
conv3_kernel[5][1][2][4]=	38236	;
conv3_kernel[5][1][3][0]=	98799	;
conv3_kernel[5][1][3][1]=	11978	;
conv3_kernel[5][1][3][2]=	-13236	;
conv3_kernel[5][1][3][3]=	24607	;
conv3_kernel[5][1][3][4]=	10127	;
conv3_kernel[5][1][4][0]=	86210	;
conv3_kernel[5][1][4][1]=	25848	;
conv3_kernel[5][1][4][2]=	19666	;
conv3_kernel[5][1][4][3]=	2068	;
conv3_kernel[5][1][4][4]=	-21561	;
conv3_kernel[6][0][0][0]=	-11692	;
conv3_kernel[6][0][0][1]=	-47628	;
conv3_kernel[6][0][0][2]=	-24463	;
conv3_kernel[6][0][0][3]=	5810	;
conv3_kernel[6][0][0][4]=	35474	;
conv3_kernel[6][0][1][0]=	-15800	;
conv3_kernel[6][0][1][1]=	17652	;
conv3_kernel[6][0][1][2]=	9209	;
conv3_kernel[6][0][1][3]=	9117	;
conv3_kernel[6][0][1][4]=	23907	;
conv3_kernel[6][0][2][0]=	17750	;
conv3_kernel[6][0][2][1]=	-1872	;
conv3_kernel[6][0][2][2]=	-14020	;
conv3_kernel[6][0][2][3]=	59833	;
conv3_kernel[6][0][2][4]=	18700	;
conv3_kernel[6][0][3][0]=	-8467	;
conv3_kernel[6][0][3][1]=	18841	;
conv3_kernel[6][0][3][2]=	-6475	;
conv3_kernel[6][0][3][3]=	24627	;
conv3_kernel[6][0][3][4]=	38623	;
conv3_kernel[6][0][4][0]=	30913	;
conv3_kernel[6][0][4][1]=	-11561	;
conv3_kernel[6][0][4][2]=	-490	;
conv3_kernel[6][0][4][3]=	8984	;
conv3_kernel[6][0][4][4]=	-9724	;
conv3_kernel[6][1][0][0]=	44584	;
conv3_kernel[6][1][0][1]=	7747	;
conv3_kernel[6][1][0][2]=	-31678	;
conv3_kernel[6][1][0][3]=	-73307	;
conv3_kernel[6][1][0][4]=	-37601	;
conv3_kernel[6][1][1][0]=	-20901	;
conv3_kernel[6][1][1][1]=	1945	;
conv3_kernel[6][1][1][2]=	-6526	;
conv3_kernel[6][1][1][3]=	-10796	;
conv3_kernel[6][1][1][4]=	-9396	;
conv3_kernel[6][1][2][0]=	40396	;
conv3_kernel[6][1][2][1]=	13680	;
conv3_kernel[6][1][2][2]=	17962	;
conv3_kernel[6][1][2][3]=	69467	;
conv3_kernel[6][1][2][4]=	10156	;
conv3_kernel[6][1][3][0]=	45961	;
conv3_kernel[6][1][3][1]=	15461	;
conv3_kernel[6][1][3][2]=	9625	;
conv3_kernel[6][1][3][3]=	22914	;
conv3_kernel[6][1][3][4]=	49763	;
conv3_kernel[6][1][4][0]=	-31808	;
conv3_kernel[6][1][4][1]=	-15741	;
conv3_kernel[6][1][4][2]=	-11754	;
conv3_kernel[6][1][4][3]=	-40347	;
conv3_kernel[6][1][4][4]=	22677	;
conv3_kernel[7][0][0][0]=	-15445	;
conv3_kernel[7][0][0][1]=	-528	;
conv3_kernel[7][0][0][2]=	-42489	;
conv3_kernel[7][0][0][3]=	-22083	;
conv3_kernel[7][0][0][4]=	-4048	;
conv3_kernel[7][0][1][0]=	-72642	;
conv3_kernel[7][0][1][1]=	4472	;
conv3_kernel[7][0][1][2]=	18527	;
conv3_kernel[7][0][1][3]=	9247	;
conv3_kernel[7][0][1][4]=	4124	;
conv3_kernel[7][0][2][0]=	13186	;
conv3_kernel[7][0][2][1]=	12738	;
conv3_kernel[7][0][2][2]=	8781	;
conv3_kernel[7][0][2][3]=	7240	;
conv3_kernel[7][0][2][4]=	16863	;
conv3_kernel[7][0][3][0]=	25172	;
conv3_kernel[7][0][3][1]=	2918	;
conv3_kernel[7][0][3][2]=	-2268	;
conv3_kernel[7][0][3][3]=	-23649	;
conv3_kernel[7][0][3][4]=	-63897	;
conv3_kernel[7][0][4][0]=	-2401	;
conv3_kernel[7][0][4][1]=	2443	;
conv3_kernel[7][0][4][2]=	-14784	;
conv3_kernel[7][0][4][3]=	6602	;
conv3_kernel[7][0][4][4]=	34102	;
conv3_kernel[7][1][0][0]=	9899	;
conv3_kernel[7][1][0][1]=	41261	;
conv3_kernel[7][1][0][2]=	5170	;
conv3_kernel[7][1][0][3]=	1762	;
conv3_kernel[7][1][0][4]=	35683	;
conv3_kernel[7][1][1][0]=	40056	;
conv3_kernel[7][1][1][1]=	4927	;
conv3_kernel[7][1][1][2]=	8680	;
conv3_kernel[7][1][1][3]=	8970	;
conv3_kernel[7][1][1][4]=	15003	;
conv3_kernel[7][1][2][0]=	-38296	;
conv3_kernel[7][1][2][1]=	-27717	;
conv3_kernel[7][1][2][2]=	34904	;
conv3_kernel[7][1][2][3]=	57065	;
conv3_kernel[7][1][2][4]=	-6587	;
conv3_kernel[7][1][3][0]=	-23637	;
conv3_kernel[7][1][3][1]=	24328	;
conv3_kernel[7][1][3][2]=	36238	;
conv3_kernel[7][1][3][3]=	22001	;
conv3_kernel[7][1][3][4]=	-43452	;
conv3_kernel[7][1][4][0]=	37628	;
conv3_kernel[7][1][4][1]=	20697	;
conv3_kernel[7][1][4][2]=	27738	;
conv3_kernel[7][1][4][3]=	-10468	;
conv3_kernel[7][1][4][4]=	-71243	;
conv3_kernel[8][0][0][0]=	-78206	;
conv3_kernel[8][0][0][1]=	-30105	;
conv3_kernel[8][0][0][2]=	15198	;
conv3_kernel[8][0][0][3]=	-3412	;
conv3_kernel[8][0][0][4]=	22703	;
conv3_kernel[8][0][1][0]=	-118736	;
conv3_kernel[8][0][1][1]=	2534	;
conv3_kernel[8][0][1][2]=	2188	;
conv3_kernel[8][0][1][3]=	4900	;
conv3_kernel[8][0][1][4]=	-8055	;
conv3_kernel[8][0][2][0]=	22848	;
conv3_kernel[8][0][2][1]=	-18457	;
conv3_kernel[8][0][2][2]=	16309	;
conv3_kernel[8][0][2][3]=	13214	;
conv3_kernel[8][0][2][4]=	41408	;
conv3_kernel[8][0][3][0]=	-2370	;
conv3_kernel[8][0][3][1]=	-3072	;
conv3_kernel[8][0][3][2]=	9908	;
conv3_kernel[8][0][3][3]=	-15808	;
conv3_kernel[8][0][3][4]=	-2881	;
conv3_kernel[8][0][4][0]=	18125	;
conv3_kernel[8][0][4][1]=	7152	;
conv3_kernel[8][0][4][2]=	-2209	;
conv3_kernel[8][0][4][3]=	7952	;
conv3_kernel[8][0][4][4]=	-5112	;
conv3_kernel[8][1][0][0]=	58717	;
conv3_kernel[8][1][0][1]=	41351	;
conv3_kernel[8][1][0][2]=	3181	;
conv3_kernel[8][1][0][3]=	-6577	;
conv3_kernel[8][1][0][4]=	31179	;
conv3_kernel[8][1][1][0]=	26011	;
conv3_kernel[8][1][1][1]=	6671	;
conv3_kernel[8][1][1][2]=	10460	;
conv3_kernel[8][1][1][3]=	27893	;
conv3_kernel[8][1][1][4]=	32165	;
conv3_kernel[8][1][2][0]=	6027	;
conv3_kernel[8][1][2][1]=	-33849	;
conv3_kernel[8][1][2][2]=	-40861	;
conv3_kernel[8][1][2][3]=	-16048	;
conv3_kernel[8][1][2][4]=	-33000	;
conv3_kernel[8][1][3][0]=	-17884	;
conv3_kernel[8][1][3][1]=	-14434	;
conv3_kernel[8][1][3][2]=	-16260	;
conv3_kernel[8][1][3][3]=	-344	;
conv3_kernel[8][1][3][4]=	-27558	;
conv3_kernel[8][1][4][0]=	-77622	;
conv3_kernel[8][1][4][1]=	9690	;
conv3_kernel[8][1][4][2]=	9122	;
conv3_kernel[8][1][4][3]=	10762	;
conv3_kernel[8][1][4][4]=	-61352	;
conv3_kernel[9][0][0][0]=	43725	;
conv3_kernel[9][0][0][1]=	-28892	;
conv3_kernel[9][0][0][2]=	-29118	;
conv3_kernel[9][0][0][3]=	-50560	;
conv3_kernel[9][0][0][4]=	-24092	;
conv3_kernel[9][0][1][0]=	41712	;
conv3_kernel[9][0][1][1]=	-18171	;
conv3_kernel[9][0][1][2]=	17308	;
conv3_kernel[9][0][1][3]=	18636	;
conv3_kernel[9][0][1][4]=	8762	;
conv3_kernel[9][0][2][0]=	-3230	;
conv3_kernel[9][0][2][1]=	-14584	;
conv3_kernel[9][0][2][2]=	71790	;
conv3_kernel[9][0][2][3]=	41731	;
conv3_kernel[9][0][2][4]=	423	;
conv3_kernel[9][0][3][0]=	-19181	;
conv3_kernel[9][0][3][1]=	-15999	;
conv3_kernel[9][0][3][2]=	43236	;
conv3_kernel[9][0][3][3]=	-30887	;
conv3_kernel[9][0][3][4]=	1057	;
conv3_kernel[9][0][4][0]=	3677	;
conv3_kernel[9][0][4][1]=	-38994	;
conv3_kernel[9][0][4][2]=	44639	;
conv3_kernel[9][0][4][3]=	24321	;
conv3_kernel[9][0][4][4]=	-22893	;
conv3_kernel[9][1][0][0]=	-7461	;
conv3_kernel[9][1][0][1]=	13288	;
conv3_kernel[9][1][0][2]=	45337	;
conv3_kernel[9][1][0][3]=	-37364	;
conv3_kernel[9][1][0][4]=	-8693	;
conv3_kernel[9][1][1][0]=	-4714	;
conv3_kernel[9][1][1][1]=	-12704	;
conv3_kernel[9][1][1][2]=	11649	;
conv3_kernel[9][1][1][3]=	-26076	;
conv3_kernel[9][1][1][4]=	-35449	;
conv3_kernel[9][1][2][0]=	-2502	;
conv3_kernel[9][1][2][1]=	-12169	;
conv3_kernel[9][1][2][2]=	29407	;
conv3_kernel[9][1][2][3]=	-3359	;
conv3_kernel[9][1][2][4]=	-1224	;
conv3_kernel[9][1][3][0]=	17362	;
conv3_kernel[9][1][3][1]=	6907	;
conv3_kernel[9][1][3][2]=	4353	;
conv3_kernel[9][1][3][3]=	3868	;
conv3_kernel[9][1][3][4]=	2836	;
conv3_kernel[9][1][4][0]=	14653	;
conv3_kernel[9][1][4][1]=	27144	;
conv3_kernel[9][1][4][2]=	1145	;
conv3_kernel[9][1][4][3]=	-3637	;
conv3_kernel[9][1][4][4]=	-13515	;
connect_matrix [0][0]=	-44394	;
connect_matrix [0][1]=	50367	;
connect_matrix [0][2]=	-6900	;
connect_matrix [0][3]=	-39843	;
connect_matrix [0][4]=	6683	;
connect_matrix [0][5]=	-7904	;
connect_matrix [0][6]=	-2725	;
connect_matrix [0][7]=	-1845	;
connect_matrix [0][8]=	25947	;
connect_matrix [0][9]=	-24563	;
connect_matrix [1][0]=	54820	;
connect_matrix [1][1]=	-18012	;
connect_matrix [1][2]=	-51769	;
connect_matrix [1][3]=	-40161	;
connect_matrix [1][4]=	-240	;
connect_matrix [1][5]=	19585	;
connect_matrix [1][6]=	20510	;
connect_matrix [1][7]=	-96414	;
connect_matrix [1][8]=	50850	;
connect_matrix [1][9]=	75383	;
connect_matrix [2][0]=	20945	;
connect_matrix [2][1]=	43469	;
connect_matrix [2][2]=	-1930	;
connect_matrix [2][3]=	18999	;
connect_matrix [2][4]=	-46407	;
connect_matrix [2][5]=	25047	;
connect_matrix [2][6]=	5853	;
connect_matrix [2][7]=	-22550	;
connect_matrix [2][8]=	-57976	;
connect_matrix [2][9]=	-2688	;
connect_matrix [3][0]=	-13977	;
connect_matrix [3][1]=	-1577	;
connect_matrix [3][2]=	-33035	;
connect_matrix [3][3]=	-543	;
connect_matrix [3][4]=	-8813	;
connect_matrix [3][5]=	48601	;
connect_matrix [3][6]=	-13513	;
connect_matrix [3][7]=	22296	;
connect_matrix [3][8]=	-46548	;
connect_matrix [3][9]=	22834	;
connect_matrix [4][0]=	-236	;
connect_matrix [4][1]=	-18743	;
connect_matrix [4][2]=	-5619	;
connect_matrix [4][3]=	-16907	;
connect_matrix [4][4]=	-34460	;
connect_matrix [4][5]=	-47534	;
connect_matrix [4][6]=	65334	;
connect_matrix [4][7]=	28847	;
connect_matrix [4][8]=	-20143	;
connect_matrix [4][9]=	23340	;
connect_matrix [5][0]=	18191	;
connect_matrix [5][1]=	-32763	;
connect_matrix [5][2]=	-34887	;
connect_matrix [5][3]=	-12803	;
connect_matrix [5][4]=	43388	;
connect_matrix [5][5]=	25155	;
connect_matrix [5][6]=	-7476	;
connect_matrix [5][7]=	20243	;
connect_matrix [5][8]=	-6480	;
connect_matrix [5][9]=	-38567	;
connect_matrix [6][0]=	-53547	;
connect_matrix [6][1]=	26538	;
connect_matrix [6][2]=	21059	;
connect_matrix [6][3]=	9517	;
connect_matrix [6][4]=	63155	;
connect_matrix [6][5]=	-93191	;
connect_matrix [6][6]=	13262	;
connect_matrix [6][7]=	-13934	;
connect_matrix [6][8]=	-14771	;
connect_matrix [6][9]=	-15990	;
connect_matrix [7][0]=	-32317	;
connect_matrix [7][1]=	-44323	;
connect_matrix [7][2]=	55377	;
connect_matrix [7][3]=	20148	;
connect_matrix [7][4]=	-5002	;
connect_matrix [7][5]=	28865	;
connect_matrix [7][6]=	-360	;
connect_matrix [7][7]=	-39861	;
connect_matrix [7][8]=	28069	;
connect_matrix [7][9]=	17126	;
connect_matrix [8][0]=	7073	;
connect_matrix [8][1]=	-2065	;
connect_matrix [8][2]=	2440	;
connect_matrix [8][3]=	58941	;
connect_matrix [8][4]=	-14024	;
connect_matrix [8][5]=	-9566	;
connect_matrix [8][6]=	-29282	;
connect_matrix [8][7]=	11909	;
connect_matrix [8][8]=	11518	;
connect_matrix [8][9]=	-9402	;
connect_matrix [9][0]=	27500	;
connect_matrix [9][1]=	-7133	;
connect_matrix [9][2]=	38437	;
connect_matrix [9][3]=	-20361	;
connect_matrix [9][4]=	-11531	;
connect_matrix [9][5]=	-23813	;
connect_matrix [9][6]=	-36144	;
connect_matrix [9][7]=	43373	;
connect_matrix [9][8]=	-32217	;
connect_matrix [9][9]=	17533	;





end
//     end
// endmodule