// module kernel_matrix_trained(conv1_kernel,conv2_kernel,conv3_kernel,connect_matrix);
//     parameter bitwidth=32;
//     output reg signed [bitwidth-1:0] conv1_kernel [1:0][4:0][4:0];
// 	output reg signed [bitwidth-1:0] conv2_kernel [1:0][1:0][4:0][4:0];
// 	output reg signed [bitwidth-1:0] conv3_kernel [9:0][1:0][4:0][4:0];
// 	output reg signed [bitwidth-1:0] connect_matrix [9:0][9:0];
//     always@(*) begin
// initial begin
assign conv1_kernel[0][0][0]=	-146	;
assign conv1_kernel[0][0][1]=	-101	;
assign conv1_kernel[0][0][2]=	46	;
assign conv1_kernel[0][0][3]=	-25	;
assign conv1_kernel[0][0][4]=	53	;
assign conv1_kernel[0][1][0]=	-180	;
assign conv1_kernel[0][1][1]=	48	;
assign conv1_kernel[0][1][2]=	45	;
assign conv1_kernel[0][1][3]=	47	;
assign conv1_kernel[0][1][4]=	25	;
assign conv1_kernel[0][2][0]=	-142	;
assign conv1_kernel[0][2][1]=	137	;
assign conv1_kernel[0][2][2]=	76	;
assign conv1_kernel[0][2][3]=	73	;
assign conv1_kernel[0][2][4]=	-10	;
assign conv1_kernel[0][3][0]=	-54	;
assign conv1_kernel[0][3][1]=	31	;
assign conv1_kernel[0][3][2]=	63	;
assign conv1_kernel[0][3][3]=	33	;
assign conv1_kernel[0][3][4]=	9	;
assign conv1_kernel[0][4][0]=	-35	;
assign conv1_kernel[0][4][1]=	68	;
assign conv1_kernel[0][4][2]=	-13	;
assign conv1_kernel[0][4][3]=	-28	;
assign conv1_kernel[0][4][4]=	-71	;
assign conv1_kernel[1][0][0]=	28	;
assign conv1_kernel[1][0][1]=	9	;
assign conv1_kernel[1][0][2]=	14	;
assign conv1_kernel[1][0][3]=	-24	;
assign conv1_kernel[1][0][4]=	-32	;
assign conv1_kernel[1][1][0]=	53	;
assign conv1_kernel[1][1][1]=	18	;
assign conv1_kernel[1][1][2]=	-4	;
assign conv1_kernel[1][1][3]=	1	;
assign conv1_kernel[1][1][4]=	-8	;
assign conv1_kernel[1][2][0]=	46	;
assign conv1_kernel[1][2][1]=	57	;
assign conv1_kernel[1][2][2]=	4	;
assign conv1_kernel[1][2][3]=	1	;
assign conv1_kernel[1][2][4]=	61	;
assign conv1_kernel[1][3][0]=	-12	;
assign conv1_kernel[1][3][1]=	84	;
assign conv1_kernel[1][3][2]=	134	;
assign conv1_kernel[1][3][3]=	56	;
assign conv1_kernel[1][3][4]=	13	;
assign conv1_kernel[1][4][0]=	-1	;
assign conv1_kernel[1][4][1]=	-11	;
assign conv1_kernel[1][4][2]=	4	;
assign conv1_kernel[1][4][3]=	30	;
assign conv1_kernel[1][4][4]=	31	;
assign conv2_kernel[0][0][0][0]=	22	;
assign conv2_kernel[0][0][0][1]=	54	;
assign conv2_kernel[0][0][0][2]=	69	;
assign conv2_kernel[0][0][0][3]=	0	;
assign conv2_kernel[0][0][0][4]=	-6	;
assign conv2_kernel[0][0][1][0]=	-70	;
assign conv2_kernel[0][0][1][1]=	50	;
assign conv2_kernel[0][0][1][2]=	35	;
assign conv2_kernel[0][0][1][3]=	-23	;
assign conv2_kernel[0][0][1][4]=	-24	;
assign conv2_kernel[0][0][2][0]=	16	;
assign conv2_kernel[0][0][2][1]=	-29	;
assign conv2_kernel[0][0][2][2]=	-10	;
assign conv2_kernel[0][0][2][3]=	6	;
assign conv2_kernel[0][0][2][4]=	45	;
assign conv2_kernel[0][0][3][0]=	28	;
assign conv2_kernel[0][0][3][1]=	5	;
assign conv2_kernel[0][0][3][2]=	-1	;
assign conv2_kernel[0][0][3][3]=	60	;
assign conv2_kernel[0][0][3][4]=	22	;
assign conv2_kernel[0][0][4][0]=	2	;
assign conv2_kernel[0][0][4][1]=	-60	;
assign conv2_kernel[0][0][4][2]=	-79	;
assign conv2_kernel[0][0][4][3]=	-114	;
assign conv2_kernel[0][0][4][4]=	-17	;
assign conv2_kernel[0][1][0][0]=	-61	;
assign conv2_kernel[0][1][0][1]=	-29	;
assign conv2_kernel[0][1][0][2]=	8	;
assign conv2_kernel[0][1][0][3]=	32	;
assign conv2_kernel[0][1][0][4]=	-55	;
assign conv2_kernel[0][1][1][0]=	-82	;
assign conv2_kernel[0][1][1][1]=	0	;
assign conv2_kernel[0][1][1][2]=	6	;
assign conv2_kernel[0][1][1][3]=	26	;
assign conv2_kernel[0][1][1][4]=	62	;
assign conv2_kernel[0][1][2][0]=	63	;
assign conv2_kernel[0][1][2][1]=	117	;
assign conv2_kernel[0][1][2][2]=	137	;
assign conv2_kernel[0][1][2][3]=	158	;
assign conv2_kernel[0][1][2][4]=	46	;
assign conv2_kernel[0][1][3][0]=	-36	;
assign conv2_kernel[0][1][3][1]=	-54	;
assign conv2_kernel[0][1][3][2]=	-1	;
assign conv2_kernel[0][1][3][3]=	-60	;
assign conv2_kernel[0][1][3][4]=	-181	;
assign conv2_kernel[0][1][4][0]=	-17	;
assign conv2_kernel[0][1][4][1]=	19	;
assign conv2_kernel[0][1][4][2]=	-58	;
assign conv2_kernel[0][1][4][3]=	-90	;
assign conv2_kernel[0][1][4][4]=	3	;
assign conv2_kernel[1][0][0][0]=	81	;
assign conv2_kernel[1][0][0][1]=	56	;
assign conv2_kernel[1][0][0][2]=	-30	;
assign conv2_kernel[1][0][0][3]=	-60	;
assign conv2_kernel[1][0][0][4]=	-24	;
assign conv2_kernel[1][0][1][0]=	-68	;
assign conv2_kernel[1][0][1][1]=	-94	;
assign conv2_kernel[1][0][1][2]=	55	;
assign conv2_kernel[1][0][1][3]=	-4	;
assign conv2_kernel[1][0][1][4]=	-58	;
assign conv2_kernel[1][0][2][0]=	-75	;
assign conv2_kernel[1][0][2][1]=	-68	;
assign conv2_kernel[1][0][2][2]=	46	;
assign conv2_kernel[1][0][2][3]=	49	;
assign conv2_kernel[1][0][2][4]=	23	;
assign conv2_kernel[1][0][3][0]=	19	;
assign conv2_kernel[1][0][3][1]=	-40	;
assign conv2_kernel[1][0][3][2]=	-123	;
assign conv2_kernel[1][0][3][3]=	-7	;
assign conv2_kernel[1][0][3][4]=	8	;
assign conv2_kernel[1][0][4][0]=	30	;
assign conv2_kernel[1][0][4][1]=	17	;
assign conv2_kernel[1][0][4][2]=	12	;
assign conv2_kernel[1][0][4][3]=	-5	;
assign conv2_kernel[1][0][4][4]=	7	;
assign conv2_kernel[1][1][0][0]=	-95	;
assign conv2_kernel[1][1][0][1]=	-64	;
assign conv2_kernel[1][1][0][2]=	-83	;
assign conv2_kernel[1][1][0][3]=	-86	;
assign conv2_kernel[1][1][0][4]=	-97	;
assign conv2_kernel[1][1][1][0]=	-23	;
assign conv2_kernel[1][1][1][1]=	-117	;
assign conv2_kernel[1][1][1][2]=	21	;
assign conv2_kernel[1][1][1][3]=	38	;
assign conv2_kernel[1][1][1][4]=	71	;
assign conv2_kernel[1][1][2][0]=	248	;
assign conv2_kernel[1][1][2][1]=	216	;
assign conv2_kernel[1][1][2][2]=	94	;
assign conv2_kernel[1][1][2][3]=	10	;
assign conv2_kernel[1][1][2][4]=	70	;
assign conv2_kernel[1][1][3][0]=	-99	;
assign conv2_kernel[1][1][3][1]=	33	;
assign conv2_kernel[1][1][3][2]=	0	;
assign conv2_kernel[1][1][3][3]=	29	;
assign conv2_kernel[1][1][3][4]=	-22	;
assign conv2_kernel[1][1][4][0]=	-146	;
assign conv2_kernel[1][1][4][1]=	-26	;
assign conv2_kernel[1][1][4][2]=	28	;
assign conv2_kernel[1][1][4][3]=	20	;
assign conv2_kernel[1][1][4][4]=	-7	;
assign conv3_kernel[0][0][0][0]=	-131	;
assign conv3_kernel[0][0][0][1]=	-30	;
assign conv3_kernel[0][0][0][2]=	38	;
assign conv3_kernel[0][0][0][3]=	49	;
assign conv3_kernel[0][0][0][4]=	11	;
assign conv3_kernel[0][0][1][0]=	-58	;
assign conv3_kernel[0][0][1][1]=	-6	;
assign conv3_kernel[0][0][1][2]=	10	;
assign conv3_kernel[0][0][1][3]=	-13	;
assign conv3_kernel[0][0][1][4]=	35	;
assign conv3_kernel[0][0][2][0]=	56	;
assign conv3_kernel[0][0][2][1]=	35	;
assign conv3_kernel[0][0][2][2]=	40	;
assign conv3_kernel[0][0][2][3]=	14	;
assign conv3_kernel[0][0][2][4]=	2	;
assign conv3_kernel[0][0][3][0]=	25	;
assign conv3_kernel[0][0][3][1]=	-9	;
assign conv3_kernel[0][0][3][2]=	63	;
assign conv3_kernel[0][0][3][3]=	-45	;
assign conv3_kernel[0][0][3][4]=	27	;
assign conv3_kernel[0][0][4][0]=	13	;
assign conv3_kernel[0][0][4][1]=	-32	;
assign conv3_kernel[0][0][4][2]=	14	;
assign conv3_kernel[0][0][4][3]=	4	;
assign conv3_kernel[0][0][4][4]=	3	;
assign conv3_kernel[0][1][0][0]=	-38	;
assign conv3_kernel[0][1][0][1]=	40	;
assign conv3_kernel[0][1][0][2]=	28	;
assign conv3_kernel[0][1][0][3]=	-71	;
assign conv3_kernel[0][1][0][4]=	-35	;
assign conv3_kernel[0][1][1][0]=	-144	;
assign conv3_kernel[0][1][1][1]=	12	;
assign conv3_kernel[0][1][1][2]=	44	;
assign conv3_kernel[0][1][1][3]=	4	;
assign conv3_kernel[0][1][1][4]=	-4	;
assign conv3_kernel[0][1][2][0]=	-96	;
assign conv3_kernel[0][1][2][1]=	-9	;
assign conv3_kernel[0][1][2][2]=	55	;
assign conv3_kernel[0][1][2][3]=	50	;
assign conv3_kernel[0][1][2][4]=	-94	;
assign conv3_kernel[0][1][3][0]=	107	;
assign conv3_kernel[0][1][3][1]=	6	;
assign conv3_kernel[0][1][3][2]=	-6	;
assign conv3_kernel[0][1][3][3]=	-33	;
assign conv3_kernel[0][1][3][4]=	49	;
assign conv3_kernel[0][1][4][0]=	164	;
assign conv3_kernel[0][1][4][1]=	-40	;
assign conv3_kernel[0][1][4][2]=	7	;
assign conv3_kernel[0][1][4][3]=	26	;
assign conv3_kernel[0][1][4][4]=	100	;
assign conv3_kernel[1][0][0][0]=	74	;
assign conv3_kernel[1][0][0][1]=	38	;
assign conv3_kernel[1][0][0][2]=	-11	;
assign conv3_kernel[1][0][0][3]=	-28	;
assign conv3_kernel[1][0][0][4]=	-165	;
assign conv3_kernel[1][0][1][0]=	25	;
assign conv3_kernel[1][0][1][1]=	24	;
assign conv3_kernel[1][0][1][2]=	-23	;
assign conv3_kernel[1][0][1][3]=	-8	;
assign conv3_kernel[1][0][1][4]=	-162	;
assign conv3_kernel[1][0][2][0]=	-100	;
assign conv3_kernel[1][0][2][1]=	-22	;
assign conv3_kernel[1][0][2][2]=	-1	;
assign conv3_kernel[1][0][2][3]=	5	;
assign conv3_kernel[1][0][2][4]=	107	;
assign conv3_kernel[1][0][3][0]=	-50	;
assign conv3_kernel[1][0][3][1]=	57	;
assign conv3_kernel[1][0][3][2]=	78	;
assign conv3_kernel[1][0][3][3]=	-2	;
assign conv3_kernel[1][0][3][4]=	83	;
assign conv3_kernel[1][0][4][0]=	78	;
assign conv3_kernel[1][0][4][1]=	75	;
assign conv3_kernel[1][0][4][2]=	-16	;
assign conv3_kernel[1][0][4][3]=	-21	;
assign conv3_kernel[1][0][4][4]=	-10	;
assign conv3_kernel[1][1][0][0]=	-52	;
assign conv3_kernel[1][1][0][1]=	-50	;
assign conv3_kernel[1][1][0][2]=	-23	;
assign conv3_kernel[1][1][0][3]=	-13	;
assign conv3_kernel[1][1][0][4]=	46	;
assign conv3_kernel[1][1][1][0]=	42	;
assign conv3_kernel[1][1][1][1]=	-12	;
assign conv3_kernel[1][1][1][2]=	-40	;
assign conv3_kernel[1][1][1][3]=	48	;
assign conv3_kernel[1][1][1][4]=	27	;
assign conv3_kernel[1][1][2][0]=	50	;
assign conv3_kernel[1][1][2][1]=	14	;
assign conv3_kernel[1][1][2][2]=	-29	;
assign conv3_kernel[1][1][2][3]=	69	;
assign conv3_kernel[1][1][2][4]=	-33	;
assign conv3_kernel[1][1][3][0]=	-70	;
assign conv3_kernel[1][1][3][1]=	52	;
assign conv3_kernel[1][1][3][2]=	-25	;
assign conv3_kernel[1][1][3][3]=	-11	;
assign conv3_kernel[1][1][3][4]=	33	;
assign conv3_kernel[1][1][4][0]=	-179	;
assign conv3_kernel[1][1][4][1]=	42	;
assign conv3_kernel[1][1][4][2]=	28	;
assign conv3_kernel[1][1][4][3]=	87	;
assign conv3_kernel[1][1][4][4]=	79	;
assign conv3_kernel[2][0][0][0]=	60	;
assign conv3_kernel[2][0][0][1]=	84	;
assign conv3_kernel[2][0][0][2]=	-32	;
assign conv3_kernel[2][0][0][3]=	35	;
assign conv3_kernel[2][0][0][4]=	-74	;
assign conv3_kernel[2][0][1][0]=	-32	;
assign conv3_kernel[2][0][1][1]=	28	;
assign conv3_kernel[2][0][1][2]=	19	;
assign conv3_kernel[2][0][1][3]=	-6	;
assign conv3_kernel[2][0][1][4]=	-86	;
assign conv3_kernel[2][0][2][0]=	15	;
assign conv3_kernel[2][0][2][1]=	15	;
assign conv3_kernel[2][0][2][2]=	-22	;
assign conv3_kernel[2][0][2][3]=	118	;
assign conv3_kernel[2][0][2][4]=	69	;
assign conv3_kernel[2][0][3][0]=	18	;
assign conv3_kernel[2][0][3][1]=	-4	;
assign conv3_kernel[2][0][3][2]=	4	;
assign conv3_kernel[2][0][3][3]=	118	;
assign conv3_kernel[2][0][3][4]=	35	;
assign conv3_kernel[2][0][4][0]=	-13	;
assign conv3_kernel[2][0][4][1]=	-43	;
assign conv3_kernel[2][0][4][2]=	-60	;
assign conv3_kernel[2][0][4][3]=	-7	;
assign conv3_kernel[2][0][4][4]=	30	;
assign conv3_kernel[2][1][0][0]=	-3	;
assign conv3_kernel[2][1][0][1]=	0	;
assign conv3_kernel[2][1][0][2]=	16	;
assign conv3_kernel[2][1][0][3]=	-1	;
assign conv3_kernel[2][1][0][4]=	30	;
assign conv3_kernel[2][1][1][0]=	58	;
assign conv3_kernel[2][1][1][1]=	20	;
assign conv3_kernel[2][1][1][2]=	22	;
assign conv3_kernel[2][1][1][3]=	58	;
assign conv3_kernel[2][1][1][4]=	19	;
assign conv3_kernel[2][1][2][0]=	-49	;
assign conv3_kernel[2][1][2][1]=	-12	;
assign conv3_kernel[2][1][2][2]=	19	;
assign conv3_kernel[2][1][2][3]=	94	;
assign conv3_kernel[2][1][2][4]=	-90	;
assign conv3_kernel[2][1][3][0]=	-14	;
assign conv3_kernel[2][1][3][1]=	13	;
assign conv3_kernel[2][1][3][2]=	30	;
assign conv3_kernel[2][1][3][3]=	-60	;
assign conv3_kernel[2][1][3][4]=	-69	;
assign conv3_kernel[2][1][4][0]=	50	;
assign conv3_kernel[2][1][4][1]=	-32	;
assign conv3_kernel[2][1][4][2]=	-68	;
assign conv3_kernel[2][1][4][3]=	-14	;
assign conv3_kernel[2][1][4][4]=	-2	;
assign conv3_kernel[3][0][0][0]=	20	;
assign conv3_kernel[3][0][0][1]=	-32	;
assign conv3_kernel[3][0][0][2]=	25	;
assign conv3_kernel[3][0][0][3]=	-27	;
assign conv3_kernel[3][0][0][4]=	-40	;
assign conv3_kernel[3][0][1][0]=	43	;
assign conv3_kernel[3][0][1][1]=	-22	;
assign conv3_kernel[3][0][1][2]=	-1	;
assign conv3_kernel[3][0][1][3]=	2	;
assign conv3_kernel[3][0][1][4]=	69	;
assign conv3_kernel[3][0][2][0]=	-1	;
assign conv3_kernel[3][0][2][1]=	-64	;
assign conv3_kernel[3][0][2][2]=	1	;
assign conv3_kernel[3][0][2][3]=	51	;
assign conv3_kernel[3][0][2][4]=	35	;
assign conv3_kernel[3][0][3][0]=	-39	;
assign conv3_kernel[3][0][3][1]=	-18	;
assign conv3_kernel[3][0][3][2]=	33	;
assign conv3_kernel[3][0][3][3]=	-117	;
assign conv3_kernel[3][0][3][4]=	-19	;
assign conv3_kernel[3][0][4][0]=	65	;
assign conv3_kernel[3][0][4][1]=	39	;
assign conv3_kernel[3][0][4][2]=	59	;
assign conv3_kernel[3][0][4][3]=	-13	;
assign conv3_kernel[3][0][4][4]=	-64	;
assign conv3_kernel[3][1][0][0]=	33	;
assign conv3_kernel[3][1][0][1]=	16	;
assign conv3_kernel[3][1][0][2]=	17	;
assign conv3_kernel[3][1][0][3]=	-81	;
assign conv3_kernel[3][1][0][4]=	34	;
assign conv3_kernel[3][1][1][0]=	-26	;
assign conv3_kernel[3][1][1][1]=	4	;
assign conv3_kernel[3][1][1][2]=	31	;
assign conv3_kernel[3][1][1][3]=	25	;
assign conv3_kernel[3][1][1][4]=	-13	;
assign conv3_kernel[3][1][2][0]=	-32	;
assign conv3_kernel[3][1][2][1]=	0	;
assign conv3_kernel[3][1][2][2]=	119	;
assign conv3_kernel[3][1][2][3]=	85	;
assign conv3_kernel[3][1][2][4]=	58	;
assign conv3_kernel[3][1][3][0]=	132	;
assign conv3_kernel[3][1][3][1]=	-16	;
assign conv3_kernel[3][1][3][2]=	-19	;
assign conv3_kernel[3][1][3][3]=	38	;
assign conv3_kernel[3][1][3][4]=	109	;
assign conv3_kernel[3][1][4][0]=	-242	;
assign conv3_kernel[3][1][4][1]=	-26	;
assign conv3_kernel[3][1][4][2]=	23	;
assign conv3_kernel[3][1][4][3]=	25	;
assign conv3_kernel[3][1][4][4]=	-23	;
assign conv3_kernel[4][0][0][0]=	-15	;
assign conv3_kernel[4][0][0][1]=	64	;
assign conv3_kernel[4][0][0][2]=	99	;
assign conv3_kernel[4][0][0][3]=	156	;
assign conv3_kernel[4][0][0][4]=	99	;
assign conv3_kernel[4][0][1][0]=	19	;
assign conv3_kernel[4][0][1][1]=	7	;
assign conv3_kernel[4][0][1][2]=	11	;
assign conv3_kernel[4][0][1][3]=	22	;
assign conv3_kernel[4][0][1][4]=	48	;
assign conv3_kernel[4][0][2][0]=	-50	;
assign conv3_kernel[4][0][2][1]=	-15	;
assign conv3_kernel[4][0][2][2]=	44	;
assign conv3_kernel[4][0][2][3]=	-71	;
assign conv3_kernel[4][0][2][4]=	-90	;
assign conv3_kernel[4][0][3][0]=	-19	;
assign conv3_kernel[4][0][3][1]=	3	;
assign conv3_kernel[4][0][3][2]=	73	;
assign conv3_kernel[4][0][3][3]=	-47	;
assign conv3_kernel[4][0][3][4]=	-2	;
assign conv3_kernel[4][0][4][0]=	17	;
assign conv3_kernel[4][0][4][1]=	-22	;
assign conv3_kernel[4][0][4][2]=	39	;
assign conv3_kernel[4][0][4][3]=	11	;
assign conv3_kernel[4][0][4][4]=	-58	;
assign conv3_kernel[4][1][0][0]=	43	;
assign conv3_kernel[4][1][0][1]=	-30	;
assign conv3_kernel[4][1][0][2]=	-68	;
assign conv3_kernel[4][1][0][3]=	-150	;
assign conv3_kernel[4][1][0][4]=	-35	;
assign conv3_kernel[4][1][1][0]=	-42	;
assign conv3_kernel[4][1][1][1]=	-27	;
assign conv3_kernel[4][1][1][2]=	-13	;
assign conv3_kernel[4][1][1][3]=	28	;
assign conv3_kernel[4][1][1][4]=	146	;
assign conv3_kernel[4][1][2][0]=	-74	;
assign conv3_kernel[4][1][2][1]=	12	;
assign conv3_kernel[4][1][2][2]=	61	;
assign conv3_kernel[4][1][2][3]=	100	;
assign conv3_kernel[4][1][2][4]=	96	;
assign conv3_kernel[4][1][3][0]=	-7	;
assign conv3_kernel[4][1][3][1]=	66	;
assign conv3_kernel[4][1][3][2]=	9	;
assign conv3_kernel[4][1][3][3]=	35	;
assign conv3_kernel[4][1][3][4]=	-20	;
assign conv3_kernel[4][1][4][0]=	-69	;
assign conv3_kernel[4][1][4][1]=	46	;
assign conv3_kernel[4][1][4][2]=	25	;
assign conv3_kernel[4][1][4][3]=	51	;
assign conv3_kernel[4][1][4][4]=	-5	;
assign conv3_kernel[5][0][0][0]=	154	;
assign conv3_kernel[5][0][0][1]=	67	;
assign conv3_kernel[5][0][0][2]=	46	;
assign conv3_kernel[5][0][0][3]=	-34	;
assign conv3_kernel[5][0][0][4]=	-67	;
assign conv3_kernel[5][0][1][0]=	89	;
assign conv3_kernel[5][0][1][1]=	23	;
assign conv3_kernel[5][0][1][2]=	7	;
assign conv3_kernel[5][0][1][3]=	-7	;
assign conv3_kernel[5][0][1][4]=	17	;
assign conv3_kernel[5][0][2][0]=	30	;
assign conv3_kernel[5][0][2][1]=	-12	;
assign conv3_kernel[5][0][2][2]=	-18	;
assign conv3_kernel[5][0][2][3]=	5	;
assign conv3_kernel[5][0][2][4]=	-45	;
assign conv3_kernel[5][0][3][0]=	0	;
assign conv3_kernel[5][0][3][1]=	26	;
assign conv3_kernel[5][0][3][2]=	-18	;
assign conv3_kernel[5][0][3][3]=	-6	;
assign conv3_kernel[5][0][3][4]=	-4	;
assign conv3_kernel[5][0][4][0]=	6	;
assign conv3_kernel[5][0][4][1]=	-47	;
assign conv3_kernel[5][0][4][2]=	-46	;
assign conv3_kernel[5][0][4][3]=	17	;
assign conv3_kernel[5][0][4][4]=	-69	;
assign conv3_kernel[5][1][0][0]=	-88	;
assign conv3_kernel[5][1][0][1]=	10	;
assign conv3_kernel[5][1][0][2]=	32	;
assign conv3_kernel[5][1][0][3]=	-6	;
assign conv3_kernel[5][1][0][4]=	12	;
assign conv3_kernel[5][1][1][0]=	-36	;
assign conv3_kernel[5][1][1][1]=	61	;
assign conv3_kernel[5][1][1][2]=	23	;
assign conv3_kernel[5][1][1][3]=	41	;
assign conv3_kernel[5][1][1][4]=	18	;
assign conv3_kernel[5][1][2][0]=	121	;
assign conv3_kernel[5][1][2][1]=	-14	;
assign conv3_kernel[5][1][2][2]=	3	;
assign conv3_kernel[5][1][2][3]=	37	;
assign conv3_kernel[5][1][2][4]=	75	;
assign conv3_kernel[5][1][3][0]=	193	;
assign conv3_kernel[5][1][3][1]=	23	;
assign conv3_kernel[5][1][3][2]=	-26	;
assign conv3_kernel[5][1][3][3]=	48	;
assign conv3_kernel[5][1][3][4]=	20	;
assign conv3_kernel[5][1][4][0]=	168	;
assign conv3_kernel[5][1][4][1]=	50	;
assign conv3_kernel[5][1][4][2]=	38	;
assign conv3_kernel[5][1][4][3]=	4	;
assign conv3_kernel[5][1][4][4]=	-42	;
assign conv3_kernel[6][0][0][0]=	-23	;
assign conv3_kernel[6][0][0][1]=	-93	;
assign conv3_kernel[6][0][0][2]=	-48	;
assign conv3_kernel[6][0][0][3]=	11	;
assign conv3_kernel[6][0][0][4]=	69	;
assign conv3_kernel[6][0][1][0]=	-31	;
assign conv3_kernel[6][0][1][1]=	34	;
assign conv3_kernel[6][0][1][2]=	18	;
assign conv3_kernel[6][0][1][3]=	18	;
assign conv3_kernel[6][0][1][4]=	47	;
assign conv3_kernel[6][0][2][0]=	35	;
assign conv3_kernel[6][0][2][1]=	-4	;
assign conv3_kernel[6][0][2][2]=	-27	;
assign conv3_kernel[6][0][2][3]=	117	;
assign conv3_kernel[6][0][2][4]=	37	;
assign conv3_kernel[6][0][3][0]=	-17	;
assign conv3_kernel[6][0][3][1]=	37	;
assign conv3_kernel[6][0][3][2]=	-13	;
assign conv3_kernel[6][0][3][3]=	48	;
assign conv3_kernel[6][0][3][4]=	75	;
assign conv3_kernel[6][0][4][0]=	60	;
assign conv3_kernel[6][0][4][1]=	-23	;
assign conv3_kernel[6][0][4][2]=	-1	;
assign conv3_kernel[6][0][4][3]=	18	;
assign conv3_kernel[6][0][4][4]=	-19	;
assign conv3_kernel[6][1][0][0]=	87	;
assign conv3_kernel[6][1][0][1]=	15	;
assign conv3_kernel[6][1][0][2]=	-62	;
assign conv3_kernel[6][1][0][3]=	-143	;
assign conv3_kernel[6][1][0][4]=	-73	;
assign conv3_kernel[6][1][1][0]=	-41	;
assign conv3_kernel[6][1][1][1]=	4	;
assign conv3_kernel[6][1][1][2]=	-13	;
assign conv3_kernel[6][1][1][3]=	-21	;
assign conv3_kernel[6][1][1][4]=	-18	;
assign conv3_kernel[6][1][2][0]=	79	;
assign conv3_kernel[6][1][2][1]=	27	;
assign conv3_kernel[6][1][2][2]=	35	;
assign conv3_kernel[6][1][2][3]=	136	;
assign conv3_kernel[6][1][2][4]=	20	;
assign conv3_kernel[6][1][3][0]=	90	;
assign conv3_kernel[6][1][3][1]=	30	;
assign conv3_kernel[6][1][3][2]=	19	;
assign conv3_kernel[6][1][3][3]=	45	;
assign conv3_kernel[6][1][3][4]=	97	;
assign conv3_kernel[6][1][4][0]=	-62	;
assign conv3_kernel[6][1][4][1]=	-31	;
assign conv3_kernel[6][1][4][2]=	-23	;
assign conv3_kernel[6][1][4][3]=	-79	;
assign conv3_kernel[6][1][4][4]=	44	;
assign conv3_kernel[7][0][0][0]=	-30	;
assign conv3_kernel[7][0][0][1]=	-1	;
assign conv3_kernel[7][0][0][2]=	-83	;
assign conv3_kernel[7][0][0][3]=	-43	;
assign conv3_kernel[7][0][0][4]=	-8	;
assign conv3_kernel[7][0][1][0]=	-142	;
assign conv3_kernel[7][0][1][1]=	9	;
assign conv3_kernel[7][0][1][2]=	36	;
assign conv3_kernel[7][0][1][3]=	18	;
assign conv3_kernel[7][0][1][4]=	8	;
assign conv3_kernel[7][0][2][0]=	26	;
assign conv3_kernel[7][0][2][1]=	25	;
assign conv3_kernel[7][0][2][2]=	17	;
assign conv3_kernel[7][0][2][3]=	14	;
assign conv3_kernel[7][0][2][4]=	33	;
assign conv3_kernel[7][0][3][0]=	49	;
assign conv3_kernel[7][0][3][1]=	6	;
assign conv3_kernel[7][0][3][2]=	-4	;
assign conv3_kernel[7][0][3][3]=	-46	;
assign conv3_kernel[7][0][3][4]=	-125	;
assign conv3_kernel[7][0][4][0]=	-5	;
assign conv3_kernel[7][0][4][1]=	5	;
assign conv3_kernel[7][0][4][2]=	-29	;
assign conv3_kernel[7][0][4][3]=	13	;
assign conv3_kernel[7][0][4][4]=	67	;
assign conv3_kernel[7][1][0][0]=	19	;
assign conv3_kernel[7][1][0][1]=	81	;
assign conv3_kernel[7][1][0][2]=	10	;
assign conv3_kernel[7][1][0][3]=	3	;
assign conv3_kernel[7][1][0][4]=	70	;
assign conv3_kernel[7][1][1][0]=	78	;
assign conv3_kernel[7][1][1][1]=	10	;
assign conv3_kernel[7][1][1][2]=	17	;
assign conv3_kernel[7][1][1][3]=	18	;
assign conv3_kernel[7][1][1][4]=	29	;
assign conv3_kernel[7][1][2][0]=	-75	;
assign conv3_kernel[7][1][2][1]=	-54	;
assign conv3_kernel[7][1][2][2]=	68	;
assign conv3_kernel[7][1][2][3]=	111	;
assign conv3_kernel[7][1][2][4]=	-13	;
assign conv3_kernel[7][1][3][0]=	-46	;
assign conv3_kernel[7][1][3][1]=	48	;
assign conv3_kernel[7][1][3][2]=	71	;
assign conv3_kernel[7][1][3][3]=	43	;
assign conv3_kernel[7][1][3][4]=	-85	;
assign conv3_kernel[7][1][4][0]=	73	;
assign conv3_kernel[7][1][4][1]=	40	;
assign conv3_kernel[7][1][4][2]=	54	;
assign conv3_kernel[7][1][4][3]=	-20	;
assign conv3_kernel[7][1][4][4]=	-139	;
assign conv3_kernel[8][0][0][0]=	-153	;
assign conv3_kernel[8][0][0][1]=	-59	;
assign conv3_kernel[8][0][0][2]=	30	;
assign conv3_kernel[8][0][0][3]=	-7	;
assign conv3_kernel[8][0][0][4]=	44	;
assign conv3_kernel[8][0][1][0]=	-232	;
assign conv3_kernel[8][0][1][1]=	5	;
assign conv3_kernel[8][0][1][2]=	4	;
assign conv3_kernel[8][0][1][3]=	10	;
assign conv3_kernel[8][0][1][4]=	-16	;
assign conv3_kernel[8][0][2][0]=	45	;
assign conv3_kernel[8][0][2][1]=	-36	;
assign conv3_kernel[8][0][2][2]=	32	;
assign conv3_kernel[8][0][2][3]=	26	;
assign conv3_kernel[8][0][2][4]=	81	;
assign conv3_kernel[8][0][3][0]=	-5	;
assign conv3_kernel[8][0][3][1]=	-6	;
assign conv3_kernel[8][0][3][2]=	19	;
assign conv3_kernel[8][0][3][3]=	-31	;
assign conv3_kernel[8][0][3][4]=	-6	;
assign conv3_kernel[8][0][4][0]=	35	;
assign conv3_kernel[8][0][4][1]=	14	;
assign conv3_kernel[8][0][4][2]=	-4	;
assign conv3_kernel[8][0][4][3]=	16	;
assign conv3_kernel[8][0][4][4]=	-10	;
assign conv3_kernel[8][1][0][0]=	115	;
assign conv3_kernel[8][1][0][1]=	81	;
assign conv3_kernel[8][1][0][2]=	6	;
assign conv3_kernel[8][1][0][3]=	-13	;
assign conv3_kernel[8][1][0][4]=	61	;
assign conv3_kernel[8][1][1][0]=	51	;
assign conv3_kernel[8][1][1][1]=	13	;
assign conv3_kernel[8][1][1][2]=	20	;
assign conv3_kernel[8][1][1][3]=	54	;
assign conv3_kernel[8][1][1][4]=	63	;
assign conv3_kernel[8][1][2][0]=	12	;
assign conv3_kernel[8][1][2][1]=	-66	;
assign conv3_kernel[8][1][2][2]=	-80	;
assign conv3_kernel[8][1][2][3]=	-31	;
assign conv3_kernel[8][1][2][4]=	-64	;
assign conv3_kernel[8][1][3][0]=	-35	;
assign conv3_kernel[8][1][3][1]=	-28	;
assign conv3_kernel[8][1][3][2]=	-32	;
assign conv3_kernel[8][1][3][3]=	-1	;
assign conv3_kernel[8][1][3][4]=	-54	;
assign conv3_kernel[8][1][4][0]=	-152	;
assign conv3_kernel[8][1][4][1]=	19	;
assign conv3_kernel[8][1][4][2]=	18	;
assign conv3_kernel[8][1][4][3]=	21	;
assign conv3_kernel[8][1][4][4]=	-120	;
assign conv3_kernel[9][0][0][0]=	85	;
assign conv3_kernel[9][0][0][1]=	-56	;
assign conv3_kernel[9][0][0][2]=	-57	;
assign conv3_kernel[9][0][0][3]=	-99	;
assign conv3_kernel[9][0][0][4]=	-47	;
assign conv3_kernel[9][0][1][0]=	81	;
assign conv3_kernel[9][0][1][1]=	-35	;
assign conv3_kernel[9][0][1][2]=	34	;
assign conv3_kernel[9][0][1][3]=	36	;
assign conv3_kernel[9][0][1][4]=	17	;
assign conv3_kernel[9][0][2][0]=	-6	;
assign conv3_kernel[9][0][2][1]=	-28	;
assign conv3_kernel[9][0][2][2]=	140	;
assign conv3_kernel[9][0][2][3]=	82	;
assign conv3_kernel[9][0][2][4]=	1	;
assign conv3_kernel[9][0][3][0]=	-37	;
assign conv3_kernel[9][0][3][1]=	-31	;
assign conv3_kernel[9][0][3][2]=	84	;
assign conv3_kernel[9][0][3][3]=	-60	;
assign conv3_kernel[9][0][3][4]=	2	;
assign conv3_kernel[9][0][4][0]=	7	;
assign conv3_kernel[9][0][4][1]=	-76	;
assign conv3_kernel[9][0][4][2]=	87	;
assign conv3_kernel[9][0][4][3]=	48	;
assign conv3_kernel[9][0][4][4]=	-45	;
assign conv3_kernel[9][1][0][0]=	-15	;
assign conv3_kernel[9][1][0][1]=	26	;
assign conv3_kernel[9][1][0][2]=	89	;
assign conv3_kernel[9][1][0][3]=	-73	;
assign conv3_kernel[9][1][0][4]=	-17	;
assign conv3_kernel[9][1][1][0]=	-9	;
assign conv3_kernel[9][1][1][1]=	-25	;
assign conv3_kernel[9][1][1][2]=	23	;
assign conv3_kernel[9][1][1][3]=	-51	;
assign conv3_kernel[9][1][1][4]=	-69	;
assign conv3_kernel[9][1][2][0]=	-5	;
assign conv3_kernel[9][1][2][1]=	-24	;
assign conv3_kernel[9][1][2][2]=	57	;
assign conv3_kernel[9][1][2][3]=	-7	;
assign conv3_kernel[9][1][2][4]=	-2	;
assign conv3_kernel[9][1][3][0]=	34	;
assign conv3_kernel[9][1][3][1]=	13	;
assign conv3_kernel[9][1][3][2]=	9	;
assign conv3_kernel[9][1][3][3]=	8	;
assign conv3_kernel[9][1][3][4]=	6	;
assign conv3_kernel[9][1][4][0]=	29	;
assign conv3_kernel[9][1][4][1]=	53	;
assign conv3_kernel[9][1][4][2]=	2	;
assign conv3_kernel[9][1][4][3]=	-7	;
assign conv3_kernel[9][1][4][4]=	-26	;
assign connect_matrix [0][0]=	-87	;
assign connect_matrix [0][1]=	98	;
assign connect_matrix [0][2]=	-13	;
assign connect_matrix [0][3]=	-78	;
assign connect_matrix [0][4]=	13	;
assign connect_matrix [0][5]=	-15	;
assign connect_matrix [0][6]=	-5	;
assign connect_matrix [0][7]=	-4	;
assign connect_matrix [0][8]=	51	;
assign connect_matrix [0][9]=	-48	;
assign connect_matrix [1][0]=	107	;
assign connect_matrix [1][1]=	-35	;
assign connect_matrix [1][2]=	-101	;
assign connect_matrix [1][3]=	-78	;
assign connect_matrix [1][4]=	0	;
assign connect_matrix [1][5]=	38	;
assign connect_matrix [1][6]=	40	;
assign connect_matrix [1][7]=	-188	;
assign connect_matrix [1][8]=	99	;
assign connect_matrix [1][9]=	147	;
assign connect_matrix [2][0]=	41	;
assign connect_matrix [2][1]=	85	;
assign connect_matrix [2][2]=	-4	;
assign connect_matrix [2][3]=	37	;
assign connect_matrix [2][4]=	-91	;
assign connect_matrix [2][5]=	49	;
assign connect_matrix [2][6]=	11	;
assign connect_matrix [2][7]=	-44	;
assign connect_matrix [2][8]=	-113	;
assign connect_matrix [2][9]=	-5	;
assign connect_matrix [3][0]=	-27	;
assign connect_matrix [3][1]=	-3	;
assign connect_matrix [3][2]=	-65	;
assign connect_matrix [3][3]=	-1	;
assign connect_matrix [3][4]=	-17	;
assign connect_matrix [3][5]=	95	;
assign connect_matrix [3][6]=	-26	;
assign connect_matrix [3][7]=	44	;
assign connect_matrix [3][8]=	-91	;
assign connect_matrix [3][9]=	45	;
assign connect_matrix [4][0]=	0	;
assign connect_matrix [4][1]=	-37	;
assign connect_matrix [4][2]=	-11	;
assign connect_matrix [4][3]=	-33	;
assign connect_matrix [4][4]=	-67	;
assign connect_matrix [4][5]=	-93	;
assign connect_matrix [4][6]=	128	;
assign connect_matrix [4][7]=	56	;
assign connect_matrix [4][8]=	-39	;
assign connect_matrix [4][9]=	46	;
assign connect_matrix [5][0]=	36	;
assign connect_matrix [5][1]=	-64	;
assign connect_matrix [5][2]=	-68	;
assign connect_matrix [5][3]=	-25	;
assign connect_matrix [5][4]=	85	;
assign connect_matrix [5][5]=	49	;
assign connect_matrix [5][6]=	-15	;
assign connect_matrix [5][7]=	40	;
assign connect_matrix [5][8]=	-13	;
assign connect_matrix [5][9]=	-75	;
assign connect_matrix [6][0]=	-105	;
assign connect_matrix [6][1]=	52	;
assign connect_matrix [6][2]=	41	;
assign connect_matrix [6][3]=	19	;
assign connect_matrix [6][4]=	123	;
assign connect_matrix [6][5]=	-182	;
assign connect_matrix [6][6]=	26	;
assign connect_matrix [6][7]=	-27	;
assign connect_matrix [6][8]=	-29	;
assign connect_matrix [6][9]=	-31	;
assign connect_matrix [7][0]=	-63	;
assign connect_matrix [7][1]=	-87	;
assign connect_matrix [7][2]=	108	;
assign connect_matrix [7][3]=	39	;
assign connect_matrix [7][4]=	-10	;
assign connect_matrix [7][5]=	56	;
assign connect_matrix [7][6]=	-1	;
assign connect_matrix [7][7]=	-78	;
assign connect_matrix [7][8]=	55	;
assign connect_matrix [7][9]=	33	;
assign connect_matrix [8][0]=	14	;
assign connect_matrix [8][1]=	-4	;
assign connect_matrix [8][2]=	5	;
assign connect_matrix [8][3]=	115	;
assign connect_matrix [8][4]=	-27	;
assign connect_matrix [8][5]=	-19	;
assign connect_matrix [8][6]=	-57	;
assign connect_matrix [8][7]=	23	;
assign connect_matrix [8][8]=	22	;
assign connect_matrix [8][9]=	-18	;
assign connect_matrix [9][0]=	54	;
assign connect_matrix [9][1]=	-14	;
assign connect_matrix [9][2]=	75	;
assign connect_matrix [9][3]=	-40	;
assign connect_matrix [9][4]=	-23	;
assign connect_matrix [9][5]=	-47	;
assign connect_matrix [9][6]=	-71	;
assign connect_matrix [9][7]=	85	;
assign connect_matrix [9][8]=	-63	;
assign connect_matrix [9][9]=	34	;




// end
//     end
// endmodule